----------------------------------------------------------------------------------
-- Company: 	ESD Group, School of Electronics, University Of Southampton
-- Engineer:	Julian A Bailey <jab@ecs.soton.ac.uk>
-- 
-- Create Date:  14th March 2011
-- Project Name: LibNeuron 2.0
-- Module Name:  Synapse Combinatorial (Com)
-- Description:  Combinatorial logic for Next State Signals in Synapse State Machine.
--
-- Dependencies: timer_com.vhd
--
-- Revision: 2.00 
--
-- Additional Comments: 14/03/2011 - Validated using testbench - JAB
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity Synapse_Com  is
  generic 
  (
     -- Module Specific Configuration Parameters
       TimerBits : natural := 32
  );
  port 
  (
     -- System Control Input Signals
       signal nReset : in std_logic;
     -- Register Inputs
        signal Reg_In : in std_logic_vector((TimerBits*2)+24 downto 0);
     -- Register Outputs  
        signal Reg_Out : out std_logic_vector((TimerBits*2)+24 downto 0);          
     -- Static Parameters
       signal Parameters  : in std_logic_vector((TimerBits*2)+15 downto 0);
     -- Combinatorial Input Signal         
       signal Axon : in std_logic;
     -- Combinatorial Output Signals
       signal SynWeightFlag : out std_logic;
       signal SynWeightOut: out std_logic_vector(15 downto 0)
  ); 
end Synapse_Com;

architecture Behavioural of Synapse_Com is
signal SynWeight   : std_logic_vector(15 downto 0);      
signal DelayTime   : std_logic_vector((TimerBits-1) downto 0);
signal DurationTime: std_logic_vector((TimerBits-1) downto 0);

signal Timer_Start : std_logic;
signal TimerPeriod : std_logic_vector((TimerBits-1) downto 0);

signal SynWeight_Q : std_logic_vector(15 downto 0);
signal LastAxon_Q  : std_logic;

constant Idle   : std_logic_vector(2 downto 0) := "001";
constant Delay  : std_logic_vector(2 downto 0) := "010";
constant Active : std_logic_vector(2 downto 0) := "100";

signal state_D : std_logic_vector(2 downto 0);
signal state_Q : std_logic_vector(2 downto 0);
signal stateprev_Q : std_logic_vector(2 downto 0);

constant Param_Synweight_Low    : natural := 0;
constant Param_SynWeight_Top    : natural := 15;
constant Param_DelayTime_Low    : natural := 16;
constant Param_DelayTime_Top    : natural := TimerBits+15;
constant Param_DurationTime_Low : natural := TimerBits+16;
constant Param_DurationTime_Top : natural := (TimerBits*2)+15;

constant Timer_Low     : natural := 0;
constant Timer_Top     : natural := (TimerBits*2)+3;
constant Finished_Pos  : natural := (TimerBits*2)+4;
constant LastAxon_Pos  : natural := (TimerBits*2)+5;
constant SynWeight_Low : natural := (TimerBits*2)+6;
constant SynWeight_Top : natural := (TimerBits*2)+21;
constant State_Low     : natural := (TimerBits*2)+22;
constant State_Top     : natural := (TimerBits*2)+24;
constant StatePrev_Low : natural := (TimerBits*2)+25;
constant StatePrev_Top : natural := (TimerBits*2)+27;

signal Finished_D : std_logic;

signal Finished_Q : std_logic;
  
begin
SynWeight    <= Parameters(Param_SynWeight_Top    downto Param_Synweight_Low);
DelayTime    <= Parameters(Param_DelayTime_Top    downto Param_DelayTime_Low);
DurationTime <= Parameters(Param_DurationTime_Top downto Param_DurationTime_Low);

Finished_Q  <= Reg_In(Finished_Pos);
LastAxon_Q  <= Reg_In(LastAxon_Pos);
SynWeight_Q <= Reg_In(SynWeight_Top downto SynWeight_Low);
State_Q     <= Reg_In(State_Top downto State_Low);
StatePrev_Q <= Reg_In(StatePrev_Top downto StatePrev_Low);

Reg_Out(Finished_Pos) <= Finished_D;
Reg_Out(LastAxon_Pos) <= Axon;
Reg_Out(SynWeight_Top downto SynWeight_Low) <= SynWeight;
Reg_Out(State_Top downto State_Low) <= State_D;
Reg_Out(StatePrev_Top downto StatePrev_Low) <= State_Q;

Timer1: entity work.Timer_Com
  generic map(TimerBits)
  port map(nReset   => nReset,
           Reg_In   => Reg_In(Timer_Top downto Timer_Low),
           Reg_Out  => Reg_Out(Timer_Top downto Timer_Low),
           Start    => Timer_Start,
           Period_In => TimerPeriod,
           Finish    => Finished_D);

OutputFlag: process(State_Q, StatePrev_Q) is
begin
  if ((State_Q = Active) AND (StatePrev_Q = Delay)) then
    SynWeightFlag <= '1';
  else
    SynWeightFlag <= '0';
  end if;
end process OutputFlag;
           
com: process (nReset, State_Q, LastAxon_Q, SynWeight_Q, Finished_Q, DelayTime, DurationTime, Axon)
begin
  if (nReset = '0') then
    Timer_Start  <= '0';
    TimerPeriod  <= (others => '0');
    SynWeightOut <= (others => '0');
    State_D <= Idle;
  else
    case State_Q is
      when Idle =>
        TimerPeriod <= DelayTime - 3;
        SynWeightOut <= (others => '0');
        Timer_Start <= '0';
        
        if ((Axon = '1') AND (LastAxon_Q = '0')) then
          State_D <= Delay;
        else
          State_D <= Idle;  
        end if;
        
      when Delay =>
        TimerPeriod <= DelayTime - 3;
        SynWeightOut <= (others => '0');
        
        if (Finished_Q = '1') then
          Timer_Start <= '0';
          State_D <= Active;
        else
          Timer_Start <= '1';
          State_D <= Delay;  
        end if;
                
      when Active =>
        TimerPeriod <= DurationTime - 3;
        SynWeightOut <= SynWeight_Q;
        
        if (Finished_Q = '1') then
          Timer_Start <= '0';
          State_D <= Idle;
        else
          Timer_Start <= '1';
          State_D <= Active;  
        end if;
                
      when others =>
        Timer_Start  <= '-';
        TimerPeriod  <= (others => '-');
        SynWeightOut <= (others => '-');
        State_D      <= (others => '-');
    end case;  
  end if;
end process com;

end architecture Behavioural;