library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

package pna_sys_pack is

-- Control Register Bits
constant RCTRL_RST  : integer := 0;
constant RCTRL_HALT : integer := 1;

end package pna_sys_pack;
