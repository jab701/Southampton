//-----------------------------------------------------------------------------
// The confidential and proprietary information contained in this file may
// only be used by a person authorised under and to the extent permitted
// by a subsisting licensing agreement from ARM Limited.
//
//            (C) COPYRIGHT 2009-2010 ARM Limited.
//                ALL RIGHTS RESERVED
//
// This entire notice must be reproduced on all copies of this file
// and copies of this file may only be made by a person if such person is
// permitted to do so under the terms of a subsisting license agreement
// from ARM Limited.
//
//      SVN Information
//
//      Checked In          : $Date:  $
//
//      Revision            : $Revision:  $
//
//      Release Information : Cortex-M0-AT510-r0p0-00rel0
//-----------------------------------------------------------------------------

//-----------------------------------------------------------------------------
// MINISWIFT CORTEX-M0 CUT-DOWN PORT-LIST AND CONFIGURATION LEVEL
// ----------------------------------------------------------------------------
//
//-----------------------------------------------------------------------------


/* Source file "MINISWIFT-rtl-mangle1.v", line 5 */
module MINISWIFT(HCLK, HRESETn, HADDR, HBURST, HMASTLOCK, HPROT, HSIZE, HTRANS, 
	HWDATA, HWRITE, HRDATA, HREADY, HRESP, NMI, IRQ, TXEV, RXEV, LOCKUP, 
	SYSRESETREQ, STCALIB, STCLKEN, SLEEPING, SLEEPDEEP, SLEEPHOLDREQn, 
	SLEEPHOLDACKn);

	output	[31:0]		HADDR;
	output	[2:0]		HBURST;
	output	[3:0]		HPROT;
	output	[2:0]		HSIZE;
	output	[1:0]		HTRANS;
	output	[31:0]		HWDATA;
	input	[31:0]		HRDATA;
	input	[3:0]		IRQ;
	input	[25:0]		STCALIB;
	input			HCLK;
	input			HRESETn;
	input			HREADY;
	input			HRESP;
	input			NMI;
	input			RXEV;
	input			STCLKEN;
	input			SLEEPHOLDREQn;
	output			HMASTLOCK;
	output			HWRITE;
	output			TXEV;
	output			LOCKUP;
	output			SYSRESETREQ;
	output			SLEEPING;
	output			SLEEPDEEP;
	output			SLEEPHOLDACKn;

	wire			In4w84;
	wire			Lo4w84;
	wire			Aq4w84;
	wire			Nr4w84;
	wire			Ws4w84;
	wire			Ju4w84;
	wire			Uv4w84;
	wire			Nx4w84;
	wire			Gz4w84;
	wire			W05w84;
	wire			P25w84;
	wire			C45w84;
	wire			V55w84;
	wire			O75w84;
	wire			H95w84;
	wire			Ab5w84;
	wire			Tc5w84;
	wire			Me5w84;
	wire			Bg5w84;
	wire			Th5w84;
	wire			Hj5w84;
	wire			Yk5w84;
	wire			Om5w84;
	wire			Eo5w84;
	wire			Up5w84;
	wire			Kr5w84;
	wire			Ct5w84;
	wire			Uu5w84;
	wire			Mw5w84;
	wire			Ey5w84;
	wire			Wz5w84;
	wire			O16w84;
	wire			G36w84;
	wire			Y46w84;
	wire			Q66w84;
	wire			I86w84;
	wire			Ba6w84;
	wire			Ub6w84;
	wire			Nd6w84;
	wire			Gf6w84;
	wire			Zg6w84;
	wire			Si6w84;
	wire			Hk6w84;
	wire			Wl6w84;
	wire			Ln6w84;
	wire			Ap6w84;
	wire			Pq6w84;
	wire			Es6w84;
	wire			Tt6w84;
	wire			Iv6w84;
	wire			Xw6w84;
	wire			My6w84;
	wire			C07w84;
	wire			S17w84;
	wire			G37w84;
	wire			Y47w84;
	wire			T67w84;
	wire			O87w84;
	wire			Ka7w84;
	wire			Fc7w84;
	wire			Ae7w84;
	wire			Vf7w84;
	wire			Qh7w84;
	wire			Lj7w84;
	wire			Gl7w84;
	wire			Bn7w84;
	wire			Wo7w84;
	wire			Rq7w84;
	wire			Ms7w84;
	wire			Iu7w84;
	wire			Ew7w84;
	wire			Ay7w84;
	wire			Wz7w84;
	wire			S18w84;
	wire			O38w84;
	wire			K58w84;
	wire			G78w84;
	wire			C98w84;
	wire			Ya8w84;
	wire			Uc8w84;
	wire			Qe8w84;
	wire			Mg8w84;
	wire			Ii8w84;
	wire			Ek8w84;
	wire			Am8w84;
	wire			Wn8w84;
	wire			Sp8w84;
	wire			Or8w84;
	wire			Kt8w84;
	wire			Gv8w84;
	wire			Cx8w84;
	wire			Xy8w84;
	wire			S09w84;
	wire			N29w84;
	wire			I49w84;
	wire			D69w84;
	wire			Y79w84;
	wire			T99w84;
	wire			Ob9w84;
	wire			Jd9w84;
	wire			Ef9w84;
	wire			Ah9w84;
	wire			Wi9w84;
	wire			Sk9w84;
	wire			Om9w84;
	wire			Ko9w84;
	wire			Gq9w84;
	wire			Cs9w84;
	wire			Yt9w84;
	wire			Uv9w84;
	wire			Qx9w84;
	wire			Mz9w84;
	wire			I1aw84;
	wire			E3aw84;
	wire			A5aw84;
	wire			W6aw84;
	wire			S8aw84;
	wire			Oaaw84;
	wire			Kcaw84;
	wire			Geaw84;
	wire			Cgaw84;
	wire			Yhaw84;
	wire			Ujaw84;
	wire			Plaw84;
	wire			Knaw84;
	wire			Fpaw84;
	wire			Araw84;
	wire			Vsaw84;
	wire			Quaw84;
	wire			Lwaw84;
	wire			Gyaw84;
	wire			B0bw84;
	wire			W1bw84;
	wire			S3bw84;
	wire			O5bw84;
	wire			K7bw84;
	wire			G9bw84;
	wire			Cbbw84;
	wire			Ycbw84;
	wire			Uebw84;
	wire			Qgbw84;
	wire			Mibw84;
	wire			Ikbw84;
	wire			Embw84;
	wire			Aobw84;
	wire			Wpbw84;
	wire			Srbw84;
	wire			Otbw84;
	wire			Kvbw84;
	wire			Gxbw84;
	wire			Czbw84;
	wire			Y0cw84;
	wire			U2cw84;
	wire			Q4cw84;
	wire			M6cw84;
	wire			H8cw84;
	wire			Cacw84;
	wire			Xbcw84;
	wire			Sdcw84;
	wire			Nfcw84;
	wire			Ihcw84;
	wire			Djcw84;
	wire			Ykcw84;
	wire			Tmcw84;
	wire			Oocw84;
	wire			Kqcw84;
	wire			Gscw84;
	wire			Cucw84;
	wire			Yvcw84;
	wire			Uxcw84;
	wire			Qzcw84;
	wire			M1dw84;
	wire			I3dw84;
	wire			E5dw84;
	wire			A7dw84;
	wire			W8dw84;
	wire			Sadw84;
	wire			Ocdw84;
	wire			Kedw84;
	wire			Ggdw84;
	wire			Cidw84;
	wire			Yjdw84;
	wire			Uldw84;
	wire			Qndw84;
	wire			Mpdw84;
	wire			Irdw84;
	wire			Etdw84;
	wire			Zudw84;
	wire			Uwdw84;
	wire			Pydw84;
	wire			K0ew84;
	wire			F2ew84;
	wire			A4ew84;
	wire			V5ew84;
	wire			Q7ew84;
	wire			L9ew84;
	wire			Gbew84;
	wire			Cdew84;
	wire			Yeew84;
	wire			Ugew84;
	wire			Qiew84;
	wire			Mkew84;
	wire			Imew84;
	wire			Eoew84;
	wire			Aqew84;
	wire			Wrew84;
	wire			Stew84;
	wire			Ovew84;
	wire			Kxew84;
	wire			Gzew84;
	wire			C1fw84;
	wire			Y2fw84;
	wire			U4fw84;
	wire			Q6fw84;
	wire			M8fw84;
	wire			Iafw84;
	wire			Ecfw84;
	wire			Aefw84;
	wire			Wffw84;
	wire			Rhfw84;
	wire			Mjfw84;
	wire			Hlfw84;
	wire			Cnfw84;
	wire			Xofw84;
	wire			Sqfw84;
	wire			Nsfw84;
	wire			Iufw84;
	wire			Dwfw84;
	wire			Yxfw84;
	wire			Uzfw84;
	wire			Q1gw84;
	wire			M3gw84;
	wire			I5gw84;
	wire			E7gw84;
	wire			A9gw84;
	wire			Wagw84;
	wire			Scgw84;
	wire			Oegw84;
	wire			Kggw84;
	wire			Gigw84;
	wire			Ckgw84;
	wire			Ylgw84;
	wire			Ungw84;
	wire			Qpgw84;
	wire			Mrgw84;
	wire			Itgw84;
	wire			Evgw84;
	wire			Axgw84;
	wire			Wygw84;
	wire			S0hw84;
	wire			O2hw84;
	wire			J4hw84;
	wire			E6hw84;
	wire			Z7hw84;
	wire			U9hw84;
	wire			Pbhw84;
	wire			Kdhw84;
	wire			Ffhw84;
	wire			Ahhw84;
	wire			Vihw84;
	wire			Qkhw84;
	wire			Mmhw84;
	wire			Iohw84;
	wire			Eqhw84;
	wire			Ashw84;
	wire			Wthw84;
	wire			Svhw84;
	wire			Oxhw84;
	wire			Kzhw84;
	wire			G1iw84;
	wire			C3iw84;
	wire			Y4iw84;
	wire			U6iw84;
	wire			Q8iw84;
	wire			Maiw84;
	wire			Iciw84;
	wire			Eeiw84;
	wire			Agiw84;
	wire			Whiw84;
	wire			Sjiw84;
	wire			Oliw84;
	wire			Kniw84;
	wire			Gpiw84;
	wire			Briw84;
	wire			Wsiw84;
	wire			Ruiw84;
	wire			Mwiw84;
	wire			Hyiw84;
	wire			C0jw84;
	wire			X1jw84;
	wire			S3jw84;
	wire			N5jw84;
	wire			I7jw84;
	wire			E9jw84;
	wire			Abjw84;
	wire			Wcjw84;
	wire			Sejw84;
	wire			Ogjw84;
	wire			Kijw84;
	wire			Gkjw84;
	wire			Cmjw84;
	wire			Ynjw84;
	wire			Upjw84;
	wire			Qrjw84;
	wire			Mtjw84;
	wire			Ivjw84;
	wire			Exjw84;
	wire			Azjw84;
	wire			W0kw84;
	wire			S2kw84;
	wire			O4kw84;
	wire			K6kw84;
	wire			G8kw84;
	wire			Cakw84;
	wire			Ybkw84;
	wire			Tdkw84;
	wire			Ofkw84;
	wire			Jhkw84;
	wire			Ejkw84;
	wire			Zkkw84;
	wire			Umkw84;
	wire			Pokw84;
	wire			Kqkw84;
	wire			Fskw84;
	wire			Aukw84;
	wire			Wvkw84;
	wire			Sxkw84;
	wire			Ozkw84;
	wire			K1lw84;
	wire			G3lw84;
	wire			C5lw84;
	wire			Y6lw84;
	wire			U8lw84;
	wire			Qalw84;
	wire			Mclw84;
	wire			Ielw84;
	wire			Eglw84;
	wire			Ailw84;
	wire			Wjlw84;
	wire			Sllw84;
	wire			Onlw84;
	wire			Kplw84;
	wire			Grlw84;
	wire			Ctlw84;
	wire			Yulw84;
	wire			Uwlw84;
	wire			Qylw84;
	wire			L0mw84;
	wire			G2mw84;
	wire			B4mw84;
	wire			W5mw84;
	wire			R7mw84;
	wire			M9mw84;
	wire			Hbmw84;
	wire			Cdmw84;
	wire			Xemw84;
	wire			Sgmw84;
	wire			Oimw84;
	wire			Kkmw84;
	wire			Gmmw84;
	wire			Comw84;
	wire			Ypmw84;
	wire			Urmw84;
	wire			Qtmw84;
	wire			Mvmw84;
	wire			Ixmw84;
	wire			Ezmw84;
	wire			A1nw84;
	wire			W2nw84;
	wire			S4nw84;
	wire			O6nw84;
	wire			K8nw84;
	wire			Ganw84;
	wire			Ccnw84;
	wire			Ydnw84;
	wire			Ufnw84;
	wire			Qhnw84;
	wire			Mjnw84;
	wire			Ilnw84;
	wire			Dnnw84;
	wire			Yonw84;
	wire			Tqnw84;
	wire			Osnw84;
	wire			Junw84;
	wire			Ewnw84;
	wire			Zxnw84;
	wire			Uznw84;
	wire			P1ow84;
	wire			K3ow84;
	wire			G5ow84;
	wire			C7ow84;
	wire			Y8ow84;
	wire			Uaow84;
	wire			Qcow84;
	wire			Meow84;
	wire			Igow84;
	wire			Eiow84;
	wire			Akow84;
	wire			Wlow84;
	wire			Snow84;
	wire			Opow84;
	wire			Krow84;
	wire			Gtow84;
	wire			Cvow84;
	wire			Ywow84;
	wire			Uyow84;
	wire			Q0pw84;
	wire			M2pw84;
	wire			I4pw84;
	wire			E6pw84;
	wire			A8pw84;
	wire			V9pw84;
	wire			Qbpw84;
	wire			Ldpw84;
	wire			Gfpw84;
	wire			Bhpw84;
	wire			Wipw84;
	wire			Rkpw84;
	wire			Mmpw84;
	wire			Hopw84;
	wire			Cqpw84;
	wire			Yrpw84;
	wire			Utpw84;
	wire			Qvpw84;
	wire			Mxpw84;
	wire			Izpw84;
	wire			E1qw84;
	wire			A3qw84;
	wire			W4qw84;
	wire			S6qw84;
	wire			O8qw84;
	wire			Kaqw84;
	wire			Gcqw84;
	wire			Ceqw84;
	wire			Yfqw84;
	wire			Uhqw84;
	wire			Qjqw84;
	wire			Mlqw84;
	wire			Inqw84;
	wire			Epqw84;
	wire			Arqw84;
	wire			Wsqw84;
	wire			Suqw84;
	wire			Nwqw84;
	wire			Iyqw84;
	wire			D0rw84;
	wire			Y1rw84;
	wire			T3rw84;
	wire			O5rw84;
	wire			J7rw84;
	wire			E9rw84;
	wire			Zarw84;
	wire			Ucrw84;
	wire			Qerw84;
	wire			Mgrw84;
	wire			Iirw84;
	wire			Ekrw84;
	wire			Amrw84;
	wire			Wnrw84;
	wire			Sprw84;
	wire			Orrw84;
	wire			Ktrw84;
	wire			Gvrw84;
	wire			Cxrw84;
	wire			Yyrw84;
	wire			U0sw84;
	wire			Q2sw84;
	wire			M4sw84;
	wire			I6sw84;
	wire			E8sw84;
	wire			Aasw84;
	wire			Wbsw84;
	wire			Sdsw84;
	wire			Ofsw84;
	wire			Khsw84;
	wire			Fjsw84;
	wire			Alsw84;
	wire			Vmsw84;
	wire			Qosw84;
	wire			Lqsw84;
	wire			Gssw84;
	wire			Busw84;
	wire			Wvsw84;
	wire			Rxsw84;
	wire			Mzsw84;
	wire			I1tw84;
	wire			E3tw84;
	wire			A5tw84;
	wire			W6tw84;
	wire			S8tw84;
	wire			Oatw84;
	wire			Kctw84;
	wire			Getw84;
	wire			Cgtw84;
	wire			Yhtw84;
	wire			Ujtw84;
	wire			Qltw84;
	wire			Mntw84;
	wire			Iptw84;
	wire			Ertw84;
	wire			Attw84;
	wire			Wutw84;
	wire			Swtw84;
	wire			Oytw84;
	wire			K0uw84;
	wire			G2uw84;
	wire			C4uw84;
	wire			X5uw84;
	wire			S7uw84;
	wire			N9uw84;
	wire			Ibuw84;
	wire			Dduw84;
	wire			Yeuw84;
	wire			Tguw84;
	wire			Oiuw84;
	wire			Jkuw84;
	wire			Emuw84;
	wire			Aouw84;
	wire			Wpuw84;
	wire			Sruw84;
	wire			Otuw84;
	wire			Kvuw84;
	wire			Gxuw84;
	wire			Czuw84;
	wire			Y0vw84;
	wire			U2vw84;
	wire			Q4vw84;
	wire			M6vw84;
	wire			I8vw84;
	wire			Eavw84;
	wire			Acvw84;
	wire			Wdvw84;
	wire			Sfvw84;
	wire			Ohvw84;
	wire			Kjvw84;
	wire			Glvw84;
	wire			Cnvw84;
	wire			Yovw84;
	wire			Uqvw84;
	wire			Psvw84;
	wire			Kuvw84;
	wire			Fwvw84;
	wire			Ayvw84;
	wire			Vzvw84;
	wire			Q1ww84;
	wire			L3ww84;
	wire			G5ww84;
	wire			B7ww84;
	wire			W8ww84;
	wire			Saww84;
	wire			Ocww84;
	wire			Keww84;
	wire			Ggww84;
	wire			Ciww84;
	wire			Yjww84;
	wire			Ulww84;
	wire			Qnww84;
	wire			Mpww84;
	wire			Irww84;
	wire			Etww84;
	wire			Avww84;
	wire			Wwww84;
	wire			Syww84;
	wire			O0xw84;
	wire			K2xw84;
	wire			G4xw84;
	wire			C6xw84;
	wire			Y7xw84;
	wire			U9xw84;
	wire			Qbxw84;
	wire			Mdxw84;
	wire			Efxw84;
	wire			Zgxw84;
	wire			Uixw84;
	wire			Pkxw84;
	wire			Kmxw84;
	wire			Foxw84;
	wire			Aqxw84;
	wire			Vrxw84;
	wire			Qtxw84;
	wire			Mvxw84;
	wire			Ixxw84;
	wire			Ezxw84;
	wire			A1yw84;
	wire			W2yw84;
	wire			S4yw84;
	wire			O6yw84;
	wire			K8yw84;
	wire			Gayw84;
	wire			Ccyw84;
	wire			Ydyw84;
	wire			Ufyw84;
	wire			Qhyw84;
	wire			Mjyw84;
	wire			Ilyw84;
	wire			Enyw84;
	wire			Apyw84;
	wire			Wqyw84;
	wire			Ssyw84;
	wire			Ouyw84;
	wire			Kwyw84;
	wire			Gyyw84;
	wire			B0zw84;
	wire			W1zw84;
	wire			R3zw84;
	wire			M5zw84;
	wire			H7zw84;
	wire			C9zw84;
	wire			Xazw84;
	wire			Sczw84;
	wire			Oezw84;
	wire			Kgzw84;
	wire			Gizw84;
	wire			Ckzw84;
	wire			Ylzw84;
	wire			Unzw84;
	wire			Qpzw84;
	wire			Mrzw84;
	wire			Itzw84;
	wire			Evzw84;
	wire			Axzw84;
	wire			Wyzw84;
	wire			S00x84;
	wire			O20x84;
	wire			K40x84;
	wire			G60x84;
	wire			C80x84;
	wire			Y90x84;
	wire			Ub0x84;
	wire			Qd0x84;
	wire			Mf0x84;
	wire			Ih0x84;
	wire			Dj0x84;
	wire			Yk0x84;
	wire			Tm0x84;
	wire			Oo0x84;
	wire			Jq0x84;
	wire			Es0x84;
	wire			Zt0x84;
	wire			Uv0x84;
	wire			Px0x84;
	wire			Kz0x84;
	wire			F11x84;
	wire			A31x84;
	wire			W41x84;
	wire			S61x84;
	wire			O81x84;
	wire			Ka1x84;
	wire			Gc1x84;
	wire			Ce1x84;
	wire			Yf1x84;
	wire			Th1x84;
	wire			Oj1x84;
	wire			Jl1x84;
	wire			En1x84;
	wire			Zo1x84;
	wire			Uq1x84;
	wire			Ps1x84;
	wire			Ku1x84;
	wire			Fw1x84;
	wire			Ay1x84;
	wire			Wz1x84;
	wire			S12x84;
	wire			O32x84;
	wire			K52x84;
	wire			G72x84;
	wire			C92x84;
	wire			Ya2x84;
	wire			Tc2x84;
	wire			Me2x84;
	wire			Ig2x84;
	wire			Bi2x84;
	wire			Uj2x84;
	wire			Ol2x84;
	wire			Fn2x84;
	wire			Zo2x84;
	wire			Tq2x84;
	wire			Ns2x84;
	wire			Hu2x84;
	wire			Bw2x84;
	wire			Vx2x84;
	wire			Pz2x84;
	wire			J13x84;
	wire			G33x84;
	wire			D53x84;
	wire			Y63x84;
	wire			R83x84;
	wire			La3x84;
	wire			Cc3x84;
	wire			Td3x84;
	wire			Kf3x84;
	wire			Bh3x84;
	wire			Yi3x84;
	wire			Vk3x84;
	wire			Qm3x84;
	wire			Oo3x84;
	wire			Mq3x84;
	wire			Js3x84;
	wire			Eu3x84;
	wire			Cw3x84;
	wire			Zx3x84;
	wire			Wz3x84;
	wire			T14x84;
	wire			Q34x84;
	wire			N54x84;
	wire			S54x84;
	wire			X54x84;
	wire			C64x84;
	wire			I64x84;
	wire			O64x84;
	wire			U64x84;
	wire			A74x84;
	wire			G74x84;
	wire			M74x84;
	wire			S74x84;
	wire			Y74x84;
	wire			E84x84;
	wire			K84x84;
	wire			Q84x84;
	wire			W84x84;
	wire			C94x84;
	wire			I94x84;
	wire			O94x84;
	wire			U94x84;
	wire			Aa4x84;
	wire			Ga4x84;
	wire			Ma4x84;
	wire			Sa4x84;
	wire			Ya4x84;
	wire			Eb4x84;
	wire			Kb4x84;
	wire			Qb4x84;
	wire			Wb4x84;
	wire			Cc4x84;
	wire			Ic4x84;
	wire			Oc4x84;
	wire			Uc4x84;
	wire			Ad4x84;
	wire			Gd4x84;
	wire			Md4x84;
	wire			Sd4x84;
	wire			Yd4x84;
	wire			Ee4x84;
	wire			Ke4x84;
	wire			Qe4x84;
	wire			We4x84;
	wire			Cf4x84;
	wire			If4x84;
	wire			Of4x84;
	wire			Uf4x84;
	wire			Ag4x84;
	wire			Gg4x84;
	wire			Mg4x84;
	wire			Sg4x84;
	wire			Yg4x84;
	wire			Eh4x84;
	wire			Kh4x84;
	wire			Qh4x84;
	wire			Wh4x84;
	wire			Ci4x84;
	wire			Ii4x84;
	wire			Oi4x84;
	wire			Ui4x84;
	wire			Aj4x84;
	wire			Gj4x84;
	wire			Mj4x84;
	wire			Sj4x84;
	wire			Yj4x84;
	wire			Ek4x84;
	wire			Kk4x84;
	wire			Qk4x84;
	wire			Wk4x84;
	wire			Cl4x84;
	wire			Il4x84;
	wire			Ol4x84;
	wire			Ul4x84;
	wire			Am4x84;
	wire			Gm4x84;
	wire			Mm4x84;
	wire			Sm4x84;
	wire			Ym4x84;
	wire			En4x84;
	wire			Kn4x84;
	wire			Qn4x84;
	wire			Wn4x84;
	wire			Co4x84;
	wire			Io4x84;
	wire			Oo4x84;
	wire			Uo4x84;
	wire			Ap4x84;
	wire			Gp4x84;
	wire			Mp4x84;
	wire			Sp4x84;
	wire			Yp4x84;
	wire			Eq4x84;
	wire			Kq4x84;
	wire			Qq4x84;
	wire			Wq4x84;
	wire			Cr4x84;
	wire			Ir4x84;
	wire			Or4x84;
	wire			Ur4x84;
	wire			As4x84;
	wire			Gs4x84;
	wire			Ms4x84;
	wire			Ss4x84;
	wire			Ys4x84;
	wire			Et4x84;
	wire			Kt4x84;
	wire			Qt4x84;
	wire			Wt4x84;
	wire			Cu4x84;
	wire			Iu4x84;
	wire			Ou4x84;
	wire			Uu4x84;
	wire			Av4x84;
	wire			Gv4x84;
	wire			Mv4x84;
	wire			Sv4x84;
	wire			Yv4x84;
	wire			Ew4x84;
	wire			Kw4x84;
	wire			Qw4x84;
	wire			Ww4x84;
	wire			Cx4x84;
	wire			Ix4x84;
	wire			Ox4x84;
	wire			Ux4x84;
	wire			Ay4x84;
	wire			Gy4x84;
	wire			My4x84;
	wire			Sy4x84;
	wire			Yy4x84;
	wire			Ez4x84;
	wire			Kz4x84;
	wire			Qz4x84;
	wire			Wz4x84;
	wire			C05x84;
	wire			I05x84;
	wire			O05x84;
	wire			U05x84;
	wire			A15x84;
	wire			G15x84;
	wire			M15x84;
	wire			S15x84;
	wire			Y15x84;
	wire			E25x84;
	wire			K25x84;
	wire			Q25x84;
	wire			W25x84;
	wire			C35x84;
	wire			I35x84;
	wire			O35x84;
	wire			U35x84;
	wire			A45x84;
	wire			G45x84;
	wire			M45x84;
	wire			S45x84;
	wire			Y45x84;
	wire			E55x84;
	wire			K55x84;
	wire			Q55x84;
	wire			W55x84;
	wire			C65x84;
	wire			I65x84;
	wire			O65x84;
	wire			U65x84;
	wire			A75x84;
	wire			G75x84;
	wire			M75x84;
	wire			S75x84;
	wire			Y75x84;
	wire			E85x84;
	wire			K85x84;
	wire			Q85x84;
	wire			W85x84;
	wire			C95x84;
	wire			I95x84;
	wire			O95x84;
	wire			U95x84;
	wire			Aa5x84;
	wire			Ga5x84;
	wire			Ma5x84;
	wire			Sa5x84;
	wire			Ya5x84;
	wire			Eb5x84;
	wire			Kb5x84;
	wire			Qb5x84;
	wire			Wb5x84;
	wire			Cc5x84;
	wire			Ic5x84;
	wire			Oc5x84;
	wire			Uc5x84;
	wire			Ad5x84;
	wire			Gd5x84;
	wire			Md5x84;
	wire			Sd5x84;
	wire			Yd5x84;
	wire			Ee5x84;
	wire			Ke5x84;
	wire			Qe5x84;
	wire			We5x84;
	wire			Cf5x84;
	wire			If5x84;
	wire			Of5x84;
	wire			Uf5x84;
	wire			Ag5x84;
	wire			Gg5x84;
	wire			Mg5x84;
	wire			Sg5x84;
	wire			Yg5x84;
	wire			Eh5x84;
	wire			Kh5x84;
	wire			Qh5x84;
	wire			Wh5x84;
	wire			Ci5x84;
	wire			Ii5x84;
	wire			Oi5x84;
	wire			Ui5x84;
	wire			Aj5x84;
	wire			Gj5x84;
	wire			Mj5x84;
	wire			Sj5x84;
	wire			Yj5x84;
	wire			Ek5x84;
	wire			Kk5x84;
	wire			Qk5x84;
	wire			Wk5x84;
	wire			Cl5x84;
	wire			Il5x84;
	wire			Ol5x84;
	wire			Ul5x84;
	wire			Am5x84;
	wire			Gm5x84;
	wire			Mm5x84;
	wire			Sm5x84;
	wire			Ym5x84;
	wire			En5x84;
	wire			Kn5x84;
	wire			Qn5x84;
	wire			Wn5x84;
	wire			Co5x84;
	wire			Io5x84;
	wire			Oo5x84;
	wire			Uo5x84;
	wire			Ap5x84;
	wire			Gp5x84;
	wire			Mp5x84;
	wire			Sp5x84;
	wire			Yp5x84;
	wire			Eq5x84;
	wire			Kq5x84;
	wire			Qq5x84;
	wire			Wq5x84;
	wire			Cr5x84;
	wire			Ir5x84;
	wire			Or5x84;
	wire			Ur5x84;
	wire			As5x84;
	wire			Gs5x84;
	wire			Ms5x84;
	wire			Ss5x84;
	wire			Ys5x84;
	wire			Et5x84;
	wire			Kt5x84;
	wire			Qt5x84;
	wire			Wt5x84;
	wire			Cu5x84;
	wire			Iu5x84;
	wire			Ou5x84;
	wire			Uu5x84;
	wire			Av5x84;
	wire			Gv5x84;
	wire			Mv5x84;
	wire			Sv5x84;
	wire			Yv5x84;
	wire			Ew5x84;
	wire			Kw5x84;
	wire			Qw5x84;
	wire			Ww5x84;
	wire			Cx5x84;
	wire			Ix5x84;
	wire			Ox5x84;
	wire			Ux5x84;
	wire			Ay5x84;
	wire			Gy5x84;
	wire			My5x84;
	wire			Sy5x84;
	wire			Yy5x84;
	wire			Ez5x84;
	wire			Kz5x84;
	wire			Qz5x84;
	wire			Wz5x84;
	wire			C06x84;
	wire			I06x84;
	wire			O06x84;
	wire			U06x84;
	wire			A16x84;
	wire			G16x84;
	wire			M16x84;
	wire			S16x84;
	wire			Y16x84;
	wire			E26x84;
	wire			K26x84;
	wire			Q26x84;
	wire			W26x84;
	wire			C36x84;
	wire			I36x84;
	wire			O36x84;
	wire			U36x84;
	wire			A46x84;
	wire			G46x84;
	wire			M46x84;
	wire			S46x84;
	wire			Y46x84;
	wire			E56x84;
	wire			K56x84;
	wire			Q56x84;
	wire			W56x84;
	wire			C66x84;
	wire			I66x84;
	wire			O66x84;
	wire			U66x84;
	wire			A76x84;
	wire			G76x84;
	wire			M76x84;
	wire			S76x84;
	wire			Y76x84;
	wire			E86x84;
	wire			K86x84;
	wire			Q86x84;
	wire			W86x84;
	wire			C96x84;
	wire			I96x84;
	wire			O96x84;
	wire			U96x84;
	wire			Aa6x84;
	wire			Ga6x84;
	wire			Ma6x84;
	wire			Sa6x84;
	wire			Ya6x84;
	wire			Eb6x84;
	wire			Kb6x84;
	wire			Qb6x84;
	wire			Wb6x84;
	wire			Cc6x84;
	wire			Ic6x84;
	wire			Oc6x84;
	wire			Uc6x84;
	wire			Ad6x84;
	wire			Gd6x84;
	wire			Md6x84;
	wire			Sd6x84;
	wire			Yd6x84;
	wire			Ee6x84;
	wire			Ke6x84;
	wire			Qe6x84;
	wire			We6x84;
	wire			Cf6x84;
	wire			If6x84;
	wire			Of6x84;
	wire			Uf6x84;
	wire			Ag6x84;
	wire			Gg6x84;
	wire			Mg6x84;
	wire			Sg6x84;
	wire			Yg6x84;
	wire			Eh6x84;
	wire			Kh6x84;
	wire			Qh6x84;
	wire			Wh6x84;
	wire			Ci6x84;
	wire			Ii6x84;
	wire			Oi6x84;
	wire			Ui6x84;
	wire			Aj6x84;
	wire			Gj6x84;
	wire			Mj6x84;
	wire			Sj6x84;
	wire			Yj6x84;
	wire			Ek6x84;
	wire			Kk6x84;
	wire			Qk6x84;
	wire			Wk6x84;
	wire			Cl6x84;
	wire			Il6x84;
	wire			Ol6x84;
	wire			Ul6x84;
	wire			Am6x84;
	wire			Gm6x84;
	wire			Mm6x84;
	wire			Sm6x84;
	wire			Ym6x84;
	wire			En6x84;
	wire			Kn6x84;
	wire			Qn6x84;
	wire			Wn6x84;
	wire			Co6x84;
	wire			Io6x84;
	wire			Oo6x84;
	wire			Uo6x84;
	wire			Ap6x84;
	wire			Gp6x84;
	wire			Mp6x84;
	wire			Sp6x84;
	wire			Yp6x84;
	wire			Eq6x84;
	wire			Kq6x84;
	wire			Qq6x84;
	wire			Wq6x84;
	wire			Cr6x84;
	wire			Ir6x84;
	wire			Or6x84;
	wire			Ur6x84;
	wire			As6x84;
	wire			Gs6x84;
	wire			Ms6x84;
	wire			Ss6x84;
	wire			Ys6x84;
	wire			Et6x84;
	wire			Kt6x84;
	wire			Qt6x84;
	wire			Wt6x84;
	wire			Cu6x84;
	wire			Iu6x84;
	wire			Ou6x84;
	wire			Uu6x84;
	wire			Av6x84;
	wire			Gv6x84;
	wire			Mv6x84;
	wire			Sv6x84;
	wire			Yv6x84;
	wire			Ew6x84;
	wire			Kw6x84;
	wire			Qw6x84;
	wire			Ww6x84;
	wire			Cx6x84;
	wire			Ix6x84;
	wire			Ox6x84;
	wire			Ux6x84;
	wire			Ay6x84;
	wire			Gy6x84;
	wire			My6x84;
	wire			Sy6x84;
	wire			Yy6x84;
	wire			Ez6x84;
	wire			Kz6x84;
	wire			Qz6x84;
	wire			Wz6x84;
	wire			C07x84;
	wire			I07x84;
	wire			O07x84;
	wire			U07x84;
	wire			A17x84;
	wire			G17x84;
	wire			M17x84;
	wire			S17x84;
	wire			Y17x84;
	wire			E27x84;
	wire			K27x84;
	wire			Q27x84;
	wire			W27x84;
	wire			C37x84;
	wire			I37x84;
	wire			O37x84;
	wire			U37x84;
	wire			A47x84;
	wire			G47x84;
	wire			M47x84;
	wire			S47x84;
	wire			Y47x84;
	wire			E57x84;
	wire			K57x84;
	wire			Q57x84;
	wire			W57x84;
	wire			C67x84;
	wire			I67x84;
	wire			O67x84;
	wire			U67x84;
	wire			A77x84;
	wire			G77x84;
	wire			M77x84;
	wire			S77x84;
	wire			Y77x84;
	wire			E87x84;
	wire			K87x84;
	wire			Q87x84;
	wire			W87x84;
	wire			C97x84;
	wire			I97x84;
	wire			O97x84;
	wire			U97x84;
	wire			Aa7x84;
	wire			Ga7x84;
	wire			Ma7x84;
	wire			Sa7x84;
	wire			Ya7x84;
	wire			Eb7x84;
	wire			Kb7x84;
	wire			Qb7x84;
	wire			Wb7x84;
	wire			Cc7x84;
	wire			Ic7x84;
	wire			Oc7x84;
	wire			Uc7x84;
	wire			Ad7x84;
	wire			Gd7x84;
	wire			Md7x84;
	wire			Sd7x84;
	wire			Yd7x84;
	wire			Ee7x84;
	wire			Ke7x84;
	wire			Qe7x84;
	wire			We7x84;
	wire			Cf7x84;
	wire			If7x84;
	wire			Of7x84;
	wire			Uf7x84;
	wire			Ag7x84;
	wire			Gg7x84;
	wire			Mg7x84;
	wire			Sg7x84;
	wire			Yg7x84;
	wire			Eh7x84;
	wire			Kh7x84;
	wire			Qh7x84;
	wire			Wh7x84;
	wire			Ci7x84;
	wire			Ii7x84;
	wire			Oi7x84;
	wire			Ui7x84;
	wire			Aj7x84;
	wire			Gj7x84;
	wire			Mj7x84;
	wire			Sj7x84;
	wire			Yj7x84;
	wire			Ek7x84;
	wire			Kk7x84;
	wire			Qk7x84;
	wire			Wk7x84;
	wire			Cl7x84;
	wire			Il7x84;
	wire			Ol7x84;
	wire			Ul7x84;
	wire			Am7x84;
	wire			Gm7x84;
	wire			Mm7x84;
	wire			Sm7x84;
	wire			Ym7x84;
	wire			En7x84;
	wire			Kn7x84;
	wire			Qn7x84;
	wire			Wn7x84;
	wire			Co7x84;
	wire			Io7x84;
	wire			Oo7x84;
	wire			Uo7x84;
	wire			Ap7x84;
	wire			Gp7x84;
	wire			Mp7x84;
	wire			Sp7x84;
	wire			Yp7x84;
	wire			Eq7x84;
	wire			Kq7x84;
	wire			Qq7x84;
	wire			Wq7x84;
	wire			Cr7x84;
	wire			Ir7x84;
	wire			Or7x84;
	wire			Ur7x84;
	wire			As7x84;
	wire			Gs7x84;
	wire			Ms7x84;
	wire			Ss7x84;
	wire			Ys7x84;
	wire			Et7x84;
	wire			Kt7x84;
	wire			Qt7x84;
	wire			Wt7x84;
	wire			Cu7x84;
	wire			Iu7x84;
	wire			Ou7x84;
	wire			Uu7x84;
	wire			Av7x84;
	wire			Gv7x84;
	wire			Mv7x84;
	wire			Sv7x84;
	wire			Yv7x84;
	wire			Ew7x84;
	wire			Kw7x84;
	wire			Qw7x84;
	wire			Ww7x84;
	wire			Cx7x84;
	wire			Ix7x84;
	wire			Ox7x84;
	wire			Ux7x84;
	wire			Ay7x84;
	wire			Gy7x84;
	wire			My7x84;
	wire			Sy7x84;
	wire			Yy7x84;
	wire			Ez7x84;
	wire			Kz7x84;
	wire			Qz7x84;
	wire			Wz7x84;
	wire			C08x84;
	wire			I08x84;
	wire			O08x84;
	wire			U08x84;
	wire			A18x84;
	wire			G18x84;
	wire			M18x84;
	wire			S18x84;
	wire			Y18x84;
	wire			E28x84;
	wire			K28x84;
	wire			Q28x84;
	wire			W28x84;
	wire			C38x84;
	wire			I38x84;
	wire			O38x84;
	wire			U38x84;
	wire			A48x84;
	wire			G48x84;
	wire			M48x84;
	wire			S48x84;
	wire			Y48x84;
	wire			E58x84;
	wire			K58x84;
	wire			Q58x84;
	wire			W58x84;
	wire			C68x84;
	wire			I68x84;
	wire			O68x84;
	wire			U68x84;
	wire			A78x84;
	wire			G78x84;
	wire			M78x84;
	wire			S78x84;
	wire			Y78x84;
	wire			E88x84;
	wire			K88x84;
	wire			Q88x84;
	wire			W88x84;
	wire			C98x84;
	wire			I98x84;
	wire			O98x84;
	wire			U98x84;
	wire			Aa8x84;
	wire			Ga8x84;
	wire			Ma8x84;
	wire			Sa8x84;
	wire			Ya8x84;
	wire			Eb8x84;
	wire			Kb8x84;
	wire			Qb8x84;
	wire			Wb8x84;
	wire			Cc8x84;
	wire			Ic8x84;
	wire			Oc8x84;
	wire			Uc8x84;
	wire			Ad8x84;
	wire			Gd8x84;
	wire			Md8x84;
	wire			Sd8x84;
	wire			Yd8x84;
	wire			Ee8x84;
	wire			Ke8x84;
	wire			Qe8x84;
	wire			We8x84;
	wire			Cf8x84;
	wire			If8x84;
	wire			Of8x84;
	wire			Uf8x84;
	wire			Ag8x84;
	wire			Gg8x84;
	wire			Mg8x84;
	wire			Sg8x84;
	wire			Yg8x84;
	wire			Eh8x84;
	wire			Kh8x84;
	wire			Qh8x84;
	wire			Wh8x84;
	wire			Ci8x84;
	wire			Ii8x84;
	wire			Oi8x84;
	wire			Ui8x84;
	wire			Aj8x84;
	wire			Gj8x84;
	wire			Mj8x84;
	wire			Sj8x84;
	wire			Yj8x84;
	wire			Ek8x84;
	wire			Kk8x84;
	wire			Qk8x84;
	wire			Wk8x84;
	wire			Cl8x84;
	wire			Il8x84;
	wire			Ol8x84;
	wire			Ul8x84;
	wire			Am8x84;
	wire			Gm8x84;
	wire			Mm8x84;
	wire			Sm8x84;
	wire			Ym8x84;
	wire			En8x84;
	wire			Kn8x84;
	wire			Qn8x84;
	wire			Wn8x84;
	wire			Co8x84;
	wire			Io8x84;
	wire			Oo8x84;
	wire			Uo8x84;
	wire			Ap8x84;
	wire			Gp8x84;
	wire			Mp8x84;
	wire			Sp8x84;
	wire			Yp8x84;
	wire			Eq8x84;
	wire			Kq8x84;
	wire			Qq8x84;
	wire			Wq8x84;
	wire			Cr8x84;
	wire			Ir8x84;
	wire			Or8x84;
	wire			Ur8x84;
	wire			As8x84;
	wire			Gs8x84;
	wire			Ms8x84;
	wire			Ss8x84;
	wire			Ys8x84;
	wire			Et8x84;
	wire			Ru8x84;
	wire			Ew8x84;
	wire			Rx8x84;
	wire			Ez8x84;
	wire			R09x84;
	wire			E29x84;
	wire			S39x84;
	wire			G59x84;
	wire			U69x84;
	wire			I89x84;
	wire			W99x84;
	wire			Kb9x84;
	wire			Xc9x84;
	wire			Le9x84;
	wire			Zf9x84;
	wire			Nh9x84;
	wire			Bj9x84;
	wire			Pk9x84;
	wire			Dm9x84;
	wire			Rn9x84;
	wire			Fp9x84;
	wire			Tq9x84;
	wire			Hs9x84;
	wire			Vt9x84;
	wire			Jv9x84;
	wire			Xw9x84;
	wire			Ly9x84;
	wire			Zz9x84;
	wire			N1ax84;
	wire			B3ax84;
	wire			P4ax84;
	wire			D6ax84;
	wire			R7ax84;
	wire			Y7ax84;
	wire			F8ax84;
	wire			M8ax84;
	wire			T8ax84;
	wire			A9ax84;
	wire			H9ax84;
	wire			O9ax84;
	wire			V9ax84;
	wire			Caax84;
	wire			Jaax84;
	wire			Qaax84;
	wire			Xaax84;
	wire			Ebax84;
	wire			Lbax84;
	wire			Sbax84;
	wire			Zbax84;
	wire			Gcax84;
	wire			Ncax84;
	wire			Ucax84;
	wire			Bdax84;
	wire			Idax84;
	wire			Pdax84;
	wire			Wdax84;
	wire			Deax84;
	wire			Keax84;
	wire			Reax84;
	wire			Yeax84;
	wire			Ffax84;
	wire			Mfax84;
	wire			Tfax84;
	wire			Agax84;
	wire			Hgax84;
	wire			Ogax84;
	wire			Vgax84;
	wire			Chax84;
	wire			Jhax84;
	wire			Qhax84;
	wire			Xhax84;
	wire			Eiax84;
	wire			Liax84;
	wire			Siax84;
	wire			Ziax84;
	wire			Gjax84;
	wire			Njax84;
	wire			Ujax84;
	wire			Bkax84;
	wire			Ikax84;
	wire			Pkax84;
	wire			Wkax84;
	wire			Dlax84;
	wire			Klax84;
	wire			Rlax84;
	wire			Ylax84;
	wire			Fmax84;
	wire			Mmax84;
	wire			Tmax84;
	wire			Anax84;
	wire			Hnax84;
	wire			Onax84;
	wire			Vnax84;
	wire			Coax84;
	wire			Joax84;
	wire			Qoax84;
	wire			Xoax84;
	wire			Epax84;
	wire			Lpax84;
	wire			Spax84;
	wire			Zpax84;
	wire			Gqax84;
	wire			Nqax84;
	wire			Uqax84;
	wire			Brax84;
	wire			Irax84;
	wire			Prax84;
	wire			Wrax84;
	wire			Dsax84;
	wire			Ksax84;
	wire			Rsax84;
	wire			Ysax84;
	wire			Ftax84;
	wire			Mtax84;
	wire			Ttax84;
	wire			Auax84;
	wire			Huax84;
	wire			Ouax84;
	wire			Vuax84;
	wire			Cvax84;
	wire			Jvax84;
	wire			Qvax84;
	wire			Xvax84;
	wire			Ewax84;
	wire			Lwax84;
	wire			Swax84;
	wire			Zwax84;
	wire			Gxax84;
	wire			Nxax84;
	wire			Uxax84;
	wire			Byax84;
	wire			Iyax84;
	wire			Pyax84;
	wire			Wyax84;
	wire			Dzax84;
	wire			Kzax84;
	wire			Rzax84;
	wire			Yzax84;
	wire			F0bx84;
	wire			M0bx84;
	wire			T0bx84;
	wire			A1bx84;
	wire			H1bx84;
	wire			O1bx84;
	wire			V1bx84;
	wire			C2bx84;
	wire			J2bx84;
	wire			Q2bx84;
	wire			X2bx84;
	wire			E3bx84;
	wire			L3bx84;
	wire			S3bx84;
	wire			Z3bx84;
	wire			G4bx84;
	wire			N4bx84;
	wire			U4bx84;
	wire			B5bx84;
	wire			I5bx84;
	wire			P5bx84;
	wire			W5bx84;
	wire			D6bx84;
	wire			K6bx84;
	wire			R6bx84;
	wire			Y6bx84;
	wire			F7bx84;
	wire			M7bx84;
	wire			T7bx84;
	wire			A8bx84;
	wire			H8bx84;
	wire			O8bx84;
	wire			V8bx84;
	wire			C9bx84;
	wire			J9bx84;
	wire			Q9bx84;
	wire			X9bx84;
	wire			Eabx84;
	wire			Labx84;
	wire			Sabx84;
	wire			Zabx84;
	wire			Gbbx84;
	wire			Nbbx84;
	wire			Ubbx84;
	wire			Bcbx84;
	wire			Icbx84;
	wire			Pcbx84;
	wire			Wcbx84;
	wire			Ddbx84;
	wire			Kdbx84;
	wire			Rdbx84;
	wire			Ydbx84;
	wire			Febx84;
	wire			Mebx84;
	wire			Tebx84;
	wire			Afbx84;
	wire			Hfbx84;
	wire			Ofbx84;
	wire			Vfbx84;
	wire			Cgbx84;
	wire			Jgbx84;
	wire			Qgbx84;
	wire			Xgbx84;
	wire			Ehbx84;
	wire			Lhbx84;
	wire			Shbx84;
	wire			Zhbx84;
	wire			Gibx84;
	wire			Nibx84;
	wire			Uibx84;
	wire			Bjbx84;
	wire			Ijbx84;
	wire			Pjbx84;
	wire			Wjbx84;
	wire			Dkbx84;
	wire			Kkbx84;
	wire			Rkbx84;
	wire			Ykbx84;
	wire			Flbx84;
	wire			Mlbx84;
	wire			Tlbx84;
	wire			Ambx84;
	wire			Hmbx84;
	wire			Ombx84;
	wire			Vmbx84;
	wire			Cnbx84;
	wire			Jnbx84;
	wire			Qnbx84;
	wire			Xnbx84;
	wire			Eobx84;
	wire			Lobx84;
	wire			Sobx84;
	wire			Zobx84;
	wire			Gpbx84;
	wire			Npbx84;
	wire			Upbx84;
	wire			Bqbx84;
	wire			Iqbx84;
	wire			Pqbx84;
	wire			Wqbx84;
	wire			Drbx84;
	wire			Krbx84;
	wire			Rrbx84;
	wire			Yrbx84;
	wire			Fsbx84;
	wire			Msbx84;
	wire			Tsbx84;
	wire			Atbx84;
	wire			Htbx84;
	wire			Otbx84;
	wire			Vtbx84;
	wire			Cubx84;
	wire			Jubx84;
	wire			Qubx84;
	wire			Xubx84;
	wire			Evbx84;
	wire			Lvbx84;
	wire			Svbx84;
	wire			Zvbx84;
	wire			Gwbx84;
	wire			Nwbx84;
	wire			Uwbx84;
	wire			Bxbx84;
	wire			Ixbx84;
	wire			Pxbx84;
	wire			Wxbx84;
	wire			Dybx84;
	wire			Kybx84;
	wire			Rybx84;
	wire			Yybx84;
	wire			Fzbx84;
	wire			Mzbx84;
	wire			Tzbx84;
	wire			A0cx84;
	wire			H0cx84;
	wire			O0cx84;
	wire			V0cx84;
	wire			C1cx84;
	wire			J1cx84;
	wire			Q1cx84;
	wire			X1cx84;
	wire			E2cx84;
	wire			L2cx84;
	wire			S2cx84;
	wire			Z2cx84;
	wire			G3cx84;
	wire			N3cx84;
	wire			U3cx84;
	wire			B4cx84;
	wire			I4cx84;
	wire			P4cx84;
	wire			W4cx84;
	wire			D5cx84;
	wire			K5cx84;
	wire			R5cx84;
	wire			Y5cx84;
	wire			F6cx84;
	wire			M6cx84;
	wire			T6cx84;
	wire			A7cx84;
	wire			H7cx84;
	wire			O7cx84;
	wire			V7cx84;
	wire			C8cx84;
	wire			J8cx84;
	wire			Q8cx84;
	wire			X8cx84;
	wire			E9cx84;
	wire			L9cx84;
	wire			S9cx84;
	wire			Z9cx84;
	wire			Gacx84;
	wire			Nacx84;
	wire			Uacx84;
	wire			Bbcx84;
	wire			Ibcx84;
	wire			Pbcx84;
	wire			Wbcx84;
	wire			Dccx84;
	wire			Kccx84;
	wire			Rccx84;
	wire			Yccx84;
	wire			Fdcx84;
	wire			Mdcx84;
	wire			Tdcx84;
	wire			Aecx84;
	wire			Hecx84;
	wire			Oecx84;
	wire			Vecx84;
	wire			Cfcx84;
	wire			Jfcx84;
	wire			Qfcx84;
	wire			Xfcx84;
	wire			Egcx84;
	wire			Lgcx84;
	wire			Sgcx84;
	wire			Zgcx84;
	wire			Ghcx84;
	wire			Nhcx84;
	wire			Uhcx84;
	wire			Bicx84;
	wire			Iicx84;
	wire			Picx84;
	wire			Wicx84;
	wire			Djcx84;
	wire			Kjcx84;
	wire			Rjcx84;
	wire			Yjcx84;
	wire			Fkcx84;
	wire			Mkcx84;
	wire			Tkcx84;
	wire			Alcx84;
	wire			Hlcx84;
	wire			Olcx84;
	wire			Vlcx84;
	wire			Cmcx84;
	wire			Jmcx84;
	wire			Qmcx84;
	wire			Xmcx84;
	wire			Encx84;
	wire			Lncx84;
	wire			Sncx84;
	wire			Zncx84;
	wire			Gocx84;
	wire			Nocx84;
	wire			Uocx84;
	wire			Bpcx84;
	wire			Ipcx84;
	wire			Ppcx84;
	wire			Wpcx84;
	wire			Dqcx84;
	wire			Kqcx84;
	wire			Rqcx84;
	wire			Yqcx84;
	wire			Frcx84;
	wire			Mrcx84;
	wire			Trcx84;
	wire			Ascx84;
	wire			Hscx84;
	wire			Oscx84;
	wire			Vscx84;
	wire			Ctcx84;
	wire			Jtcx84;
	wire			Qtcx84;
	wire			Xtcx84;
	wire			Eucx84;
	wire			Lucx84;
	wire			Sucx84;
	wire			Zucx84;
	wire			Gvcx84;
	wire			Nvcx84;
	wire			Uvcx84;
	wire			Bwcx84;
	wire			Iwcx84;
	wire			Pwcx84;
	wire			Wwcx84;
	wire			Dxcx84;
	wire			Kxcx84;
	wire			Rxcx84;
	wire			Yxcx84;
	wire			Fycx84;
	wire			Mycx84;
	wire			Tycx84;
	wire			Azcx84;
	wire			Hzcx84;
	wire			Ozcx84;
	wire			Vzcx84;
	wire			C0dx84;
	wire			J0dx84;
	wire			Q0dx84;
	wire			X0dx84;
	wire			E1dx84;
	wire			L1dx84;
	wire			S1dx84;
	wire			Z1dx84;
	wire			G2dx84;
	wire			N2dx84;
	wire			U2dx84;
	wire			B3dx84;
	wire			I3dx84;
	wire			P3dx84;
	wire			W3dx84;
	wire			D4dx84;
	wire			K4dx84;
	wire			R4dx84;
	wire			Y4dx84;
	wire			F5dx84;
	wire			M5dx84;
	wire			T5dx84;
	wire			A6dx84;
	wire			H6dx84;
	wire			O6dx84;
	wire			V6dx84;
	wire			C7dx84;
	wire			J7dx84;
	wire			Q7dx84;
	wire			X7dx84;
	wire			E8dx84;
	wire			L8dx84;
	wire			S8dx84;
	wire			Z8dx84;
	wire			G9dx84;
	wire			N9dx84;
	wire			U9dx84;
	wire			Badx84;
	wire			Iadx84;
	wire			Padx84;
	wire			Wadx84;
	wire			Dbdx84;
	wire			Kbdx84;
	wire			Rbdx84;
	wire			Ybdx84;
	wire			Fcdx84;
	wire			Mcdx84;
	wire			Tcdx84;
	wire			Addx84;
	wire			Hddx84;
	wire			Oddx84;
	wire			Vddx84;
	wire			Cedx84;
	wire			Jedx84;
	wire			Qedx84;
	wire			Xedx84;
	wire			Efdx84;
	wire			Lfdx84;
	wire			Sfdx84;
	wire			Zfdx84;
	wire			Ggdx84;
	wire			Ngdx84;
	wire			Ugdx84;
	wire			Bhdx84;
	wire			Ihdx84;
	wire			Phdx84;
	wire			Whdx84;
	wire			Didx84;
	wire			Kidx84;
	wire			Ridx84;
	wire			Yidx84;
	wire			Fjdx84;
	wire			Mjdx84;
	wire			Tjdx84;
	wire			Akdx84;
	wire			Hkdx84;
	wire			Okdx84;
	wire			Vkdx84;
	wire			Cldx84;
	wire			Jldx84;
	wire			Qldx84;
	wire			Xldx84;
	wire			Emdx84;
	wire			Lmdx84;
	wire			Smdx84;
	wire			Zmdx84;
	wire			Gndx84;
	wire			Nndx84;
	wire			Undx84;
	wire			Bodx84;
	wire			Iodx84;
	wire			Podx84;
	wire			Wodx84;
	wire			Dpdx84;
	wire			Kpdx84;
	wire			Rpdx84;
	wire			Ypdx84;
	wire			Fqdx84;
	wire			Mqdx84;
	wire			Tqdx84;
	wire			Ardx84;
	wire			Hrdx84;
	wire			Ordx84;
	wire			Vrdx84;
	wire			Csdx84;
	wire			Jsdx84;
	wire			Qsdx84;
	wire			Xsdx84;
	wire			Etdx84;
	wire			Ltdx84;
	wire			Stdx84;
	wire			Ztdx84;
	wire			Gudx84;
	wire			Nudx84;
	wire			Uudx84;
	wire			Bvdx84;
	wire			Ivdx84;
	wire			Pvdx84;
	wire			Wvdx84;
	wire			Dwdx84;
	wire			Kwdx84;
	wire			Rwdx84;
	wire			Ywdx84;
	wire			Fxdx84;
	wire			Mxdx84;
	wire			Txdx84;
	wire			Aydx84;
	wire			Hydx84;
	wire			Oydx84;
	wire			Vydx84;
	wire			Czdx84;
	wire			Jzdx84;
	wire			Qzdx84;
	wire			Xzdx84;
	wire			E0ex84;
	wire			L0ex84;
	wire			S0ex84;
	wire			Z0ex84;
	wire			G1ex84;
	wire			N1ex84;
	wire			U1ex84;
	wire			B2ex84;
	wire			I2ex84;
	wire			P2ex84;
	wire			W2ex84;
	wire			D3ex84;
	wire			K3ex84;
	wire			R3ex84;
	wire			Y3ex84;
	wire			F4ex84;
	wire			M4ex84;
	wire			T4ex84;
	wire			A5ex84;
	wire			H5ex84;
	wire			O5ex84;
	wire			V5ex84;
	wire			C6ex84;
	wire			J6ex84;
	wire			Q6ex84;
	wire			X6ex84;
	wire			E7ex84;
	wire			L7ex84;
	wire			S7ex84;
	wire			Z7ex84;
	wire			G8ex84;
	wire			N8ex84;
	wire			U8ex84;
	wire			B9ex84;
	wire			I9ex84;
	wire			P9ex84;
	wire			W9ex84;
	wire			Daex84;
	wire			Kaex84;
	wire			Raex84;
	wire			Yaex84;
	wire			Fbex84;
	wire			Mbex84;
	wire			Tbex84;
	wire			Acex84;
	wire			Hcex84;
	wire			Ocex84;
	wire			Vcex84;
	wire			Cdex84;
	wire			Jdex84;
	wire			Qdex84;
	wire			Xdex84;
	wire			Eeex84;
	wire			Leex84;
	wire			Seex84;
	wire			Zeex84;
	wire			Gfex84;
	wire			Nfex84;
	wire			Ufex84;
	wire			Bgex84;
	wire			Igex84;
	wire			Pgex84;
	wire			Wgex84;
	wire			Dhex84;
	wire			Khex84;
	wire			Rhex84;
	wire			Yhex84;
	wire			Fiex84;
	wire			Miex84;
	wire			Tiex84;
	wire			Ajex84;
	wire			Hjex84;
	wire			Ojex84;
	wire			Vjex84;
	wire			Ckex84;
	wire			Jkex84;
	wire			Qkex84;
	wire			Xkex84;
	wire			Elex84;
	wire			Llex84;
	wire			Slex84;
	wire			Zlex84;
	wire			Gmex84;
	wire			Nmex84;
	wire			Umex84;
	wire			Bnex84;
	wire			Inex84;
	wire			Pnex84;
	wire			Wnex84;
	wire			Doex84;
	wire			Koex84;
	wire			Roex84;
	wire			Yoex84;
	wire			Fpex84;
	wire			Mpex84;
	wire			Tpex84;
	wire			Aqex84;
	wire			Hqex84;
	wire			Oqex84;
	wire			Vqex84;
	wire			Crex84;
	wire			Jrex84;
	wire			Qrex84;
	wire			Xrex84;
	wire			Esex84;
	wire			Lsex84;
	wire			Ssex84;
	wire			Zsex84;
	wire			Gtex84;
	wire			Ntex84;
	wire			Utex84;
	wire			Buex84;
	wire			Iuex84;
	wire			Puex84;
	wire			Wuex84;
	wire			Dvex84;
	wire			Kvex84;
	wire			Rvex84;
	wire			Yvex84;
	wire			Fwex84;
	wire			Mwex84;
	wire			Twex84;
	wire			Axex84;
	wire			Hxex84;
	wire			Oxex84;
	wire			Vxex84;
	wire			Cyex84;
	wire			Jyex84;
	wire			Qyex84;
	wire			Xyex84;
	wire			Ezex84;
	wire			Lzex84;
	wire			Szex84;
	wire			Zzex84;
	wire			G0fx84;
	wire			N0fx84;
	wire			U0fx84;
	wire			B1fx84;
	wire			I1fx84;
	wire			P1fx84;
	wire			W1fx84;
	wire			D2fx84;
	wire			K2fx84;
	wire			R2fx84;
	wire			Y2fx84;
	wire			F3fx84;
	wire			M3fx84;
	wire			T3fx84;
	wire			A4fx84;
	wire			H4fx84;
	wire			O4fx84;
	wire			V4fx84;
	wire			C5fx84;
	wire			J5fx84;
	wire			Q5fx84;
	wire			X5fx84;
	wire			E6fx84;
	wire			L6fx84;
	wire			S6fx84;
	wire			Z6fx84;
	wire			G7fx84;
	wire			N7fx84;
	wire			U7fx84;
	wire			B8fx84;
	wire			I8fx84;
	wire			P8fx84;
	wire			W8fx84;
	wire			D9fx84;
	wire			K9fx84;
	wire			R9fx84;
	wire			Y9fx84;
	wire			Fafx84;
	wire			Mafx84;
	wire			Tafx84;
	wire			Abfx84;
	wire			Hbfx84;
	wire			Obfx84;
	wire			Vbfx84;
	wire			Ccfx84;
	wire			Jcfx84;
	wire			Qcfx84;
	wire			Xcfx84;
	wire			Edfx84;
	wire			Ldfx84;
	wire			Sdfx84;
	wire			Zdfx84;
	wire			Gefx84;
	wire			Nefx84;
	wire			Uefx84;
	wire			Bffx84;
	wire			Iffx84;
	wire			Pffx84;
	wire			Wffx84;
	wire			Dgfx84;
	wire			Kgfx84;
	wire			Rgfx84;
	wire			Ygfx84;
	wire			Fhfx84;
	wire			Mhfx84;
	wire			Thfx84;
	wire			Aifx84;
	wire			Hifx84;
	wire			Oifx84;
	wire			Vifx84;
	wire			Cjfx84;
	wire			Jjfx84;
	wire			Qjfx84;
	wire			Xjfx84;
	wire			Ekfx84;
	wire			Lkfx84;
	wire			Skfx84;
	wire			Zkfx84;
	wire			Glfx84;
	wire			Nlfx84;
	wire			Ulfx84;
	wire			Bmfx84;
	wire			Imfx84;
	wire			Pmfx84;
	wire			Wmfx84;
	wire			Dnfx84;
	wire			Knfx84;
	wire			Rnfx84;
	wire			Ynfx84;
	wire			Fofx84;
	wire			Mofx84;
	wire			Tofx84;
	wire			Apfx84;
	wire			Hpfx84;
	wire			Opfx84;
	wire			Vpfx84;
	wire			Cqfx84;
	wire			Jqfx84;
	wire			Qqfx84;
	wire			Xqfx84;
	wire			Erfx84;
	wire			Lrfx84;
	wire			Srfx84;
	wire			Zrfx84;
	wire			Gsfx84;
	wire			Nsfx84;
	wire			Usfx84;
	wire			Btfx84;
	wire			Itfx84;
	wire			Ptfx84;
	wire			Wtfx84;
	wire			Dufx84;
	wire			Kufx84;
	wire			Rufx84;
	wire			Yufx84;
	wire			Fvfx84;
	wire			Mvfx84;
	wire			Tvfx84;
	wire			Awfx84;
	wire			Hwfx84;
	wire			Owfx84;
	wire			Vwfx84;
	wire			Cxfx84;
	wire			Jxfx84;
	wire			Qxfx84;
	wire			Xxfx84;
	wire			Eyfx84;
	wire			Lyfx84;
	wire			Syfx84;
	wire			Zyfx84;
	wire			Gzfx84;
	wire			Nzfx84;
	wire			Uzfx84;
	wire			B0gx84;
	wire			I0gx84;
	wire			P0gx84;
	wire			W0gx84;
	wire			D1gx84;
	wire			K1gx84;
	wire			R1gx84;
	wire			Y1gx84;
	wire			F2gx84;
	wire			M2gx84;
	wire			T2gx84;
	wire			A3gx84;
	wire			H3gx84;
	wire			O3gx84;
	wire			V3gx84;
	wire			C4gx84;
	wire			J4gx84;
	wire			Q4gx84;
	wire			X4gx84;
	wire			E5gx84;
	wire			L5gx84;
	wire			S5gx84;
	wire			Z5gx84;
	wire			G6gx84;
	wire			N6gx84;
	wire			U6gx84;
	wire			B7gx84;
	wire			I7gx84;
	wire			P7gx84;
	wire			W7gx84;
	wire			D8gx84;
	wire			K8gx84;
	wire			R8gx84;
	wire			Y8gx84;
	wire			F9gx84;
	wire			M9gx84;
	wire			T9gx84;
	wire			Aagx84;
	wire			Hagx84;
	wire			Oagx84;
	wire			Vagx84;
	wire			Cbgx84;
	wire			Jbgx84;
	wire			Qbgx84;
	wire			Xbgx84;
	wire			Ecgx84;
	wire			Lcgx84;
	wire			Scgx84;
	wire			Zcgx84;
	wire			Gdgx84;
	wire			Ndgx84;
	wire			Udgx84;
	wire			Begx84;
	wire			Iegx84;
	wire			Pegx84;
	wire			Wegx84;
	wire			Dfgx84;
	wire			Kfgx84;
	wire			Rfgx84;
	wire			Yfgx84;
	wire			Fggx84;
	wire			Mggx84;
	wire			Tggx84;
	wire			Ahgx84;
	wire			Hhgx84;
	wire			Ohgx84;
	wire			Vhgx84;
	wire			Cigx84;
	wire			Jigx84;
	wire			Qigx84;
	wire			Xigx84;
	wire			Ejgx84;
	wire			Ljgx84;
	wire			Sjgx84;
	wire			Zjgx84;
	wire			Gkgx84;
	wire			Nkgx84;
	wire			Ukgx84;
	wire			Blgx84;
	wire			Ilgx84;
	wire			Plgx84;
	wire			Wlgx84;
	wire			Dmgx84;
	wire			Kmgx84;
	wire			Rmgx84;
	wire			Ymgx84;
	wire			Fngx84;
	wire			Mngx84;
	wire			Tngx84;
	wire			Aogx84;
	wire			Hogx84;
	wire			Oogx84;
	wire			Vogx84;
	wire			Cpgx84;
	wire			Jpgx84;
	wire			Qpgx84;
	wire			Xpgx84;
	wire			Eqgx84;
	wire			Lqgx84;
	wire			Sqgx84;
	wire			Zqgx84;
	wire			Grgx84;
	wire			Nrgx84;
	wire			Urgx84;
	wire			Bsgx84;
	wire			Isgx84;
	wire			Psgx84;
	wire			Wsgx84;
	wire			Dtgx84;
	wire			Ktgx84;
	wire			Rtgx84;
	wire			Ytgx84;
	wire			Fugx84;
	wire			Mugx84;
	wire			Tugx84;
	wire			Avgx84;
	wire			Hvgx84;
	wire			Ovgx84;
	wire			Vvgx84;
	wire			Cwgx84;
	wire			Jwgx84;
	wire			Qwgx84;
	wire			Xwgx84;
	wire			Exgx84;
	wire			Lxgx84;
	wire			Sxgx84;
	wire			Zxgx84;
	wire			Gygx84;
	wire			Nygx84;
	wire			Uygx84;
	wire			Bzgx84;
	wire			Izgx84;
	wire			Pzgx84;
	wire			Wzgx84;
	wire			D0hx84;
	wire			K0hx84;
	wire			R0hx84;
	wire			Y0hx84;
	wire			F1hx84;
	wire			M1hx84;
	wire			T1hx84;
	wire			A2hx84;
	wire			H2hx84;
	wire			O2hx84;
	wire			V2hx84;
	wire			C3hx84;
	wire			J3hx84;
	wire			Q3hx84;
	wire			X3hx84;
	wire			E4hx84;
	wire			L4hx84;
	wire			S4hx84;
	wire			Z4hx84;
	wire			G5hx84;
	wire			N5hx84;
	wire			U5hx84;
	wire			B6hx84;
	wire			I6hx84;
	wire			P6hx84;
	wire			W6hx84;
	wire			D7hx84;
	wire			K7hx84;
	wire			R7hx84;
	wire			Y7hx84;
	wire			F8hx84;
	wire			M8hx84;
	wire			T8hx84;
	wire			A9hx84;
	wire			H9hx84;
	wire			O9hx84;
	wire			V9hx84;
	wire			Cahx84;
	wire			Jahx84;
	wire			Qahx84;
	wire			Xahx84;
	wire			Ebhx84;
	wire			Lbhx84;
	wire			Sbhx84;
	wire			Zbhx84;
	wire			Gchx84;
	wire			Nchx84;
	wire			Uchx84;
	wire			Bdhx84;
	wire			Idhx84;
	wire			Pdhx84;
	wire			Wdhx84;
	wire			Dehx84;
	wire			Kehx84;
	wire			Rehx84;
	wire			Yehx84;
	wire			Ffhx84;
	wire			Mfhx84;
	wire			Tfhx84;
	wire			Aghx84;
	wire			Hghx84;
	wire			Oghx84;
	wire			Vghx84;
	wire			Chhx84;
	wire			Jhhx84;
	wire			Qhhx84;
	wire			Xhhx84;
	wire			Eihx84;
	wire			Lihx84;
	wire			Sihx84;
	wire			Zihx84;
	wire			Gjhx84;
	wire			Njhx84;
	wire			Ujhx84;
	wire			Bkhx84;
	wire			Ikhx84;
	wire			Pkhx84;
	wire			Wkhx84;
	wire			Dlhx84;
	wire			Klhx84;
	wire			Rlhx84;
	wire			Ylhx84;
	wire			Fmhx84;
	wire			Mmhx84;
	wire			Tmhx84;
	wire			Anhx84;
	wire			Hnhx84;
	wire			Onhx84;
	wire			Vnhx84;
	wire			Cohx84;
	wire			Johx84;
	wire			Qohx84;
	wire			Xohx84;
	wire			Ephx84;
	wire			Lphx84;
	wire			Sphx84;
	wire			Zphx84;
	wire			Gqhx84;
	wire			Nqhx84;
	wire			Uqhx84;
	wire			Brhx84;
	wire			Irhx84;
	wire			Prhx84;
	wire			Wrhx84;
	wire			Dshx84;
	wire			Kshx84;
	wire			Rshx84;
	wire			Yshx84;
	wire			Fthx84;
	wire			Mthx84;
	wire			Tthx84;
	wire			Auhx84;
	wire			Huhx84;
	wire			Ouhx84;
	wire			Vuhx84;
	wire			Cvhx84;
	wire			Jvhx84;
	wire			Qvhx84;
	wire			Xvhx84;
	wire			Ewhx84;
	wire			Lwhx84;
	wire			Swhx84;
	wire			Zwhx84;
	wire			Gxhx84;
	wire			Nxhx84;
	wire			Uxhx84;
	wire			Byhx84;
	wire			Iyhx84;
	wire			Pyhx84;
	wire			Wyhx84;
	wire			Dzhx84;
	wire			Kzhx84;
	wire			Rzhx84;
	wire			Yzhx84;
	wire			F0ix84;
	wire			M0ix84;
	wire			T0ix84;
	wire			A1ix84;
	wire			H1ix84;
	wire			O1ix84;
	wire			V1ix84;
	wire			C2ix84;
	wire			J2ix84;
	wire			Q2ix84;
	wire			X2ix84;
	wire			E3ix84;
	wire			L3ix84;
	wire			S3ix84;
	wire			Z3ix84;
	wire			G4ix84;
	wire			N4ix84;
	wire			U4ix84;
	wire			B5ix84;
	wire			I5ix84;
	wire			P5ix84;
	wire			W5ix84;
	wire			D6ix84;
	wire			K6ix84;
	wire			R6ix84;
	wire			Y6ix84;
	wire			F7ix84;
	wire			M7ix84;
	wire			T7ix84;
	wire			A8ix84;
	wire			H8ix84;
	wire			O8ix84;
	wire			V8ix84;
	wire			C9ix84;
	wire			J9ix84;
	wire			Q9ix84;
	wire			X9ix84;
	wire			Eaix84;
	wire			Laix84;
	wire			Saix84;
	wire			Zaix84;
	wire			Gbix84;
	wire			Nbix84;
	wire			Ubix84;
	wire			Bcix84;
	wire			Icix84;
	wire			Pcix84;
	wire			Wcix84;
	wire			Ddix84;
	wire			Kdix84;
	wire			Rdix84;
	wire			Ydix84;
	wire			Feix84;
	wire			Meix84;
	wire			Teix84;
	wire			Afix84;
	wire			Hfix84;
	wire			Ofix84;
	wire			Vfix84;
	wire			Cgix84;
	wire			Jgix84;
	wire			Qgix84;
	wire			Xgix84;
	wire			Ehix84;
	wire			Lhix84;
	wire			Shix84;
	wire			Zhix84;
	wire			Giix84;
	wire			Niix84;
	wire			Uiix84;
	wire			Bjix84;
	wire			Ijix84;
	wire			Pjix84;
	wire			Wjix84;
	wire			Dkix84;
	wire			Kkix84;
	wire			Rkix84;
	wire			Ykix84;
	wire			Flix84;
	wire			Mlix84;
	wire			Tlix84;
	wire			Amix84;
	wire			Hmix84;
	wire			Omix84;
	wire			Vmix84;
	wire			Cnix84;
	wire			Jnix84;
	wire			Qnix84;
	wire			Xnix84;
	wire			Eoix84;
	wire			Loix84;
	wire			Soix84;
	wire			Zoix84;
	wire			Gpix84;
	wire			Npix84;
	wire			Upix84;
	wire			Bqix84;
	wire			Iqix84;
	wire			Pqix84;
	wire			Wqix84;
	wire			Drix84;
	wire			Krix84;
	wire			Rrix84;
	wire			Yrix84;
	wire			Fsix84;
	wire			Msix84;
	wire			Tsix84;
	wire			Atix84;
	wire			Htix84;
	wire			Otix84;
	wire			Vtix84;
	wire			Cuix84;
	wire			Juix84;
	wire			Quix84;
	wire			Xuix84;
	wire			Evix84;
	wire			Lvix84;
	wire			Svix84;
	wire			Zvix84;
	wire			Gwix84;
	wire			Nwix84;
	wire			Uwix84;
	wire			Bxix84;
	wire			Ixix84;
	wire			Pxix84;
	wire			Wxix84;
	wire			Dyix84;
	wire			Kyix84;
	wire			Ryix84;
	wire			Yyix84;
	wire			Fzix84;
	wire			Mzix84;
	wire			Tzix84;
	wire			A0jx84;
	wire			H0jx84;
	wire			O0jx84;
	wire			V0jx84;
	wire			C1jx84;
	wire			J1jx84;
	wire			Q1jx84;
	wire			X1jx84;
	wire			E2jx84;
	wire			L2jx84;
	wire			S2jx84;
	wire			Z2jx84;
	wire			G3jx84;
	wire			N3jx84;
	wire			U3jx84;
	wire			B4jx84;
	wire			I4jx84;
	wire			P4jx84;
	wire			W4jx84;
	wire			D5jx84;
	wire			K5jx84;
	wire			R5jx84;
	wire			Y5jx84;
	wire			F6jx84;
	wire			M6jx84;
	wire			T6jx84;
	wire			A7jx84;
	wire			H7jx84;
	wire			O7jx84;
	wire			V7jx84;
	wire			C8jx84;
	wire			J8jx84;
	wire			Q8jx84;
	wire			X8jx84;
	wire			E9jx84;
	wire			L9jx84;
	wire			S9jx84;
	wire			Z9jx84;
	wire			Gajx84;
	wire			Najx84;
	wire			Uajx84;
	wire			Bbjx84;
	wire			Ibjx84;
	wire			Pbjx84;
	wire			Wbjx84;
	wire			Dcjx84;
	wire			Kcjx84;
	wire			Rcjx84;
	wire			Ycjx84;
	wire			Fdjx84;
	wire			Mdjx84;
	wire			Tdjx84;
	wire			Aejx84;
	wire			Hejx84;
	wire			Oejx84;
	wire			Vejx84;
	wire			Cfjx84;
	wire			Jfjx84;
	wire			Qfjx84;
	wire			Xfjx84;
	wire			Egjx84;
	wire			Lgjx84;
	wire			Sgjx84;
	wire			Zgjx84;
	wire			Ghjx84;
	wire			Nhjx84;
	wire			Uhjx84;
	wire			Bijx84;
	wire			Iijx84;
	wire			Pijx84;
	wire			Wijx84;
	wire			Djjx84;
	wire			Kjjx84;
	wire			Rjjx84;
	wire			Yjjx84;
	wire			Fkjx84;
	wire			Mkjx84;
	wire			Tkjx84;
	wire			Aljx84;
	wire			Hljx84;
	wire			Oljx84;
	wire			Vljx84;
	wire			Cmjx84;
	wire			Jmjx84;
	wire			Qmjx84;
	wire			Xmjx84;
	wire			Enjx84;
	wire			Lnjx84;
	wire			Snjx84;
	wire			Znjx84;
	wire			Gojx84;
	wire			Nojx84;
	wire			Uojx84;
	wire			Bpjx84;
	wire			Ipjx84;
	wire			Ppjx84;
	wire			Wpjx84;
	wire			Dqjx84;
	wire			Kqjx84;
	wire			Rqjx84;
	wire			Yqjx84;
	wire			Frjx84;
	wire			Mrjx84;
	wire			Trjx84;
	wire			Asjx84;
	wire			Hsjx84;
	wire			Osjx84;
	wire			Vsjx84;
	wire			Ctjx84;
	wire			Jtjx84;
	wire			Qtjx84;
	wire			Xtjx84;
	wire			Eujx84;
	wire			Lujx84;
	wire			Sujx84;
	wire			Zujx84;
	wire			Gvjx84;
	wire			Nvjx84;
	wire			Uvjx84;
	wire			Bwjx84;
	wire			Iwjx84;
	wire			Pwjx84;
	wire			Wwjx84;
	wire			Dxjx84;
	wire			Kxjx84;
	wire			Rxjx84;
	wire			Yxjx84;
	wire			Fyjx84;
	wire			Myjx84;
	wire			Tyjx84;
	wire			Azjx84;
	wire			Hzjx84;
	wire			Ozjx84;
	wire			Vzjx84;
	wire			C0kx84;
	wire			J0kx84;
	wire			Q0kx84;
	wire			X0kx84;
	wire			E1kx84;
	wire			L1kx84;
	wire			S1kx84;
	wire			Z1kx84;
	wire			G2kx84;
	wire			N2kx84;
	wire			U2kx84;
	wire			B3kx84;
	wire			I3kx84;
	wire			P3kx84;
	wire			W3kx84;
	wire			D4kx84;
	wire			K4kx84;
	wire			R4kx84;
	wire			Y4kx84;
	wire			F5kx84;
	wire			M5kx84;
	wire			T5kx84;
	wire			A6kx84;
	wire			H6kx84;
	wire			O6kx84;
	wire			V6kx84;
	wire			C7kx84;
	wire			J7kx84;
	wire			Q7kx84;
	wire			X7kx84;
	wire			E8kx84;
	wire			L8kx84;
	wire			S8kx84;
	wire			Z8kx84;
	wire			G9kx84;
	wire			N9kx84;
	wire			U9kx84;
	wire			Bakx84;
	wire			Iakx84;
	wire			Pakx84;
	wire			Wakx84;
	wire			Dbkx84;
	wire			Kbkx84;
	wire			Rbkx84;
	wire			Ybkx84;
	wire			Fckx84;
	wire			Mckx84;
	wire			Tckx84;
	wire			Adkx84;
	wire			Hdkx84;
	wire			Odkx84;
	wire			Vdkx84;
	wire			Cekx84;
	wire			Jekx84;
	wire			Qekx84;
	wire			Xekx84;
	wire			Efkx84;
	wire			Lfkx84;
	wire			Sfkx84;
	wire			Zfkx84;
	wire			Ggkx84;
	wire			Ngkx84;
	wire			Ugkx84;
	wire			Bhkx84;
	wire			Ihkx84;
	wire			Phkx84;
	wire			Whkx84;
	wire			Dikx84;
	wire			Kikx84;
	wire			Rikx84;
	wire			Yikx84;
	wire			Fjkx84;
	wire			Mjkx84;
	wire			Tjkx84;
	wire			Akkx84;
	wire			Hkkx84;
	wire			Okkx84;
	wire			Vkkx84;
	wire			Clkx84;
	wire			Jlkx84;
	wire			Qlkx84;
	wire			Xlkx84;
	wire			Emkx84;
	wire			Lmkx84;
	wire			Smkx84;
	wire			Zmkx84;
	wire			Gnkx84;
	wire			Nnkx84;
	wire			Unkx84;
	wire			Bokx84;
	wire			Iokx84;
	wire			Pokx84;
	wire			Wokx84;
	wire			Dpkx84;
	wire			Kpkx84;
	wire			Rpkx84;
	wire			Ypkx84;
	wire			Fqkx84;
	wire			Mqkx84;
	wire			Tqkx84;
	wire			Arkx84;
	wire			Hrkx84;
	wire			Orkx84;
	wire			Vrkx84;
	wire			Cskx84;
	wire			Jskx84;
	wire			Qskx84;
	wire			Xskx84;
	wire			Etkx84;
	wire			Ltkx84;
	wire			Stkx84;
	wire			Ztkx84;
	wire			Gukx84;
	wire			Nukx84;
	wire			Uukx84;
	wire			Bvkx84;
	wire			Ivkx84;
	wire			Pvkx84;
	wire			Wvkx84;
	wire			Dwkx84;
	wire			Kwkx84;
	wire			Rwkx84;
	wire			Ywkx84;
	wire			Fxkx84;
	wire			Mxkx84;
	wire			Txkx84;
	wire			Aykx84;
	wire			Hykx84;
	wire			Oykx84;
	wire			Vykx84;
	wire			Czkx84;
	wire			Jzkx84;
	wire			Qzkx84;
	wire			Xzkx84;
	wire			E0lx84;
	wire			L0lx84;
	wire			S0lx84;
	wire			Z0lx84;
	wire			G1lx84;
	wire			N1lx84;
	wire			U1lx84;
	wire			B2lx84;
	wire			I2lx84;
	wire			P2lx84;
	wire			W2lx84;
	wire			D3lx84;
	wire			K3lx84;
	wire			R3lx84;
	wire			Y3lx84;
	wire			F4lx84;
	wire			M4lx84;
	wire			T4lx84;
	wire			A5lx84;
	wire			H5lx84;
	wire			O5lx84;
	wire			V5lx84;
	wire			C6lx84;
	wire			J6lx84;
	wire			Q6lx84;
	wire			X6lx84;
	wire			E7lx84;
	wire			L7lx84;
	wire			S7lx84;
	wire			Z7lx84;
	wire			G8lx84;
	wire			N8lx84;
	wire			U8lx84;
	wire			B9lx84;
	wire			I9lx84;
	wire			P9lx84;
	wire			W9lx84;
	wire			Dalx84;
	wire			Kalx84;
	wire			Ralx84;
	wire			Yalx84;
	wire			Fblx84;
	wire			Mblx84;
	wire			Tblx84;
	wire			Aclx84;
	wire			Hclx84;
	wire			Oclx84;
	wire			Vclx84;
	wire			Cdlx84;
	wire			Jdlx84;
	wire			Qdlx84;
	wire			Xdlx84;
	wire			Eelx84;
	wire			Lelx84;
	wire			Selx84;
	wire			Zelx84;
	wire			Gflx84;
	wire			Nflx84;
	wire			Uflx84;
	wire			Bglx84;
	wire			Iglx84;
	wire			Pglx84;
	wire			Wglx84;
	wire			Dhlx84;
	wire			Khlx84;
	wire			Rhlx84;
	wire			Yhlx84;
	wire			Filx84;
	wire			Milx84;
	wire			Tilx84;
	wire			Ajlx84;
	wire			Hjlx84;
	wire			Ojlx84;
	wire			Vjlx84;
	wire			Cklx84;
	wire			Jklx84;
	wire			Qklx84;
	wire			Xklx84;
	wire			Ellx84;
	wire			Lllx84;
	wire			Sllx84;
	wire			Zllx84;
	wire			Gmlx84;
	wire			Nmlx84;
	wire			Umlx84;
	wire			Bnlx84;
	wire			Inlx84;
	wire			Pnlx84;
	wire			Wnlx84;
	wire			Dolx84;
	wire			Kolx84;
	wire			Rolx84;
	wire			Yolx84;
	wire			Fplx84;
	wire			Mplx84;
	wire			Tplx84;
	wire			Aqlx84;
	wire			Hqlx84;
	wire			Oqlx84;
	wire			Vqlx84;
	wire			Crlx84;
	wire			Jrlx84;
	wire			Qrlx84;
	wire			Xrlx84;
	wire			Eslx84;
	wire			Lslx84;
	wire			Sslx84;
	wire			Zslx84;
	wire			Gtlx84;
	wire			Ntlx84;
	wire			Utlx84;
	wire			Bulx84;
	wire			Iulx84;
	wire			Pulx84;
	wire			Wulx84;
	wire			Dvlx84;
	wire			Kvlx84;
	wire			Rvlx84;
	wire			Yvlx84;
	wire			Fwlx84;
	wire			Mwlx84;
	wire			Twlx84;
	wire			Axlx84;
	wire			Hxlx84;
	wire			Oxlx84;
	wire			Vxlx84;
	wire			Cylx84;
	wire			Jylx84;
	wire			Qylx84;
	wire			Xylx84;
	wire			Ezlx84;
	wire			Lzlx84;
	wire			Szlx84;
	wire			Zzlx84;
	wire			G0mx84;
	wire			N0mx84;
	wire			U0mx84;
	wire			B1mx84;
	wire			I1mx84;
	wire			P1mx84;
	wire			W1mx84;
	wire			D2mx84;
	wire			K2mx84;
	wire			R2mx84;
	wire			Y2mx84;
	wire			F3mx84;
	wire			M3mx84;
	wire			T3mx84;
	wire			A4mx84;
	wire			H4mx84;
	wire			O4mx84;
	wire			V4mx84;
	wire			C5mx84;
	wire			J5mx84;
	wire			Q5mx84;
	wire			X5mx84;
	wire			E6mx84;
	wire			L6mx84;
	wire			S6mx84;
	wire			Z6mx84;
	wire			G7mx84;
	wire			N7mx84;
	wire			U7mx84;
	wire			B8mx84;
	wire			I8mx84;
	wire			P8mx84;
	wire			W8mx84;
	wire			D9mx84;
	wire			K9mx84;
	wire			R9mx84;
	wire			Y9mx84;
	wire			Famx84;
	wire			Mamx84;
	wire			Tamx84;
	wire			Abmx84;
	wire			Hbmx84;
	wire			Obmx84;
	wire			Vbmx84;
	wire			Ccmx84;
	wire			Jcmx84;
	wire			Qcmx84;
	wire			Xcmx84;
	wire			Edmx84;
	wire			Ldmx84;
	wire			Sdmx84;
	wire			Zdmx84;
	wire			Gemx84;
	wire			Nemx84;
	wire			Uemx84;
	wire			Bfmx84;
	wire			Ifmx84;
	wire			Pfmx84;
	wire			Wfmx84;
	wire			Dgmx84;
	wire			Kgmx84;
	wire			Rgmx84;
	wire			Ygmx84;
	wire			Fhmx84;
	wire			Mhmx84;
	wire			Thmx84;
	wire			Aimx84;
	wire			Himx84;
	wire			Oimx84;
	wire			Vimx84;
	wire			Cjmx84;
	wire			Jjmx84;
	wire			Qjmx84;
	wire			Xjmx84;
	wire			Ekmx84;
	wire			Lkmx84;
	wire			Skmx84;
	wire			Zkmx84;
	wire			Glmx84;
	wire			Nlmx84;
	wire			Ulmx84;
	wire			Bmmx84;
	wire			Immx84;
	wire			Pmmx84;
	wire			Wmmx84;
	wire			Dnmx84;
	wire			Knmx84;
	wire			Rnmx84;
	wire			Ynmx84;
	wire			Fomx84;
	wire			Momx84;
	wire			Tomx84;
	wire			Apmx84;
	wire			Hpmx84;
	wire			Opmx84;
	wire			Vpmx84;
	wire			Cqmx84;
	wire			Jqmx84;
	wire			Qqmx84;
	wire			Xqmx84;
	wire			Ermx84;
	wire			Lrmx84;
	wire			Srmx84;
	wire			Zrmx84;
	wire			Gsmx84;
	wire			Nsmx84;
	wire			Usmx84;
	wire			Btmx84;
	wire			Itmx84;
	wire			Ptmx84;
	wire			Wtmx84;
	wire			Dumx84;
	wire			Kumx84;
	wire			Rumx84;
	wire			Yumx84;
	wire			Fvmx84;
	wire			Mvmx84;
	wire			Tvmx84;
	wire			Awmx84;
	wire			Hwmx84;
	wire			Owmx84;
	wire			Vwmx84;
	wire			Cxmx84;
	wire			Jxmx84;
	wire			Qxmx84;
	wire			Xxmx84;
	wire			Eymx84;
	wire			Lymx84;
	wire			Symx84;
	wire			Zymx84;
	wire			Gzmx84;
	wire			Nzmx84;
	wire			Uzmx84;
	wire			B0nx84;
	wire			I0nx84;
	wire			P0nx84;
	wire			W0nx84;
	wire			D1nx84;
	wire			K1nx84;
	wire			R1nx84;
	wire			Y1nx84;
	wire			F2nx84;
	wire			M2nx84;
	wire			T2nx84;
	wire			A3nx84;
	wire			H3nx84;
	wire			O3nx84;
	wire			V3nx84;
	wire			C4nx84;
	wire			J4nx84;
	wire			Q4nx84;
	wire			X4nx84;
	wire			E5nx84;
	wire			L5nx84;
	wire			S5nx84;
	wire			Z5nx84;
	wire			G6nx84;
	wire			N6nx84;
	wire			U6nx84;
	wire			B7nx84;
	wire			I7nx84;
	wire			P7nx84;
	wire			W7nx84;
	wire			D8nx84;
	wire			K8nx84;
	wire			R8nx84;
	wire			Y8nx84;
	wire			F9nx84;
	wire			M9nx84;
	wire			T9nx84;
	wire			Aanx84;
	wire			Hanx84;
	wire			Oanx84;
	wire			Vanx84;
	wire			Cbnx84;
	wire			Jbnx84;
	wire			Qbnx84;
	wire			Xbnx84;
	wire			Ecnx84;
	wire			Lcnx84;
	wire			Scnx84;
	wire			Zcnx84;
	wire			Gdnx84;
	wire			Ndnx84;
	wire			Udnx84;
	wire			Benx84;
	wire			Ienx84;
	wire			Penx84;
	wire			Wenx84;
	wire			Dfnx84;
	wire			Kfnx84;
	wire			Rfnx84;
	wire			Yfnx84;
	wire			Fgnx84;
	wire			Mgnx84;
	wire			Tgnx84;
	wire			Ahnx84;
	wire			Hhnx84;
	wire			Ohnx84;
	wire			Vhnx84;
	wire			Cinx84;
	wire			Jinx84;
	wire			Qinx84;
	wire			Xinx84;
	wire			Ejnx84;
	wire			Ljnx84;
	wire			Sjnx84;
	wire			Zjnx84;
	wire			Gknx84;
	wire			Nknx84;
	wire			Uknx84;
	wire			Blnx84;
	wire			Ilnx84;
	wire			Plnx84;
	wire			Wlnx84;
	wire			Dmnx84;
	wire			Kmnx84;
	wire			Rmnx84;
	wire			Ymnx84;
	wire			Fnnx84;
	wire			Mnnx84;
	wire			Tnnx84;
	wire			Aonx84;
	wire			Honx84;
	wire			Oonx84;
	wire			Vonx84;
	wire			Cpnx84;
	wire			Jpnx84;
	wire			Qpnx84;
	wire			Xpnx84;
	wire			Eqnx84;
	wire			Lqnx84;
	wire			Sqnx84;
	wire			Zqnx84;
	wire			Grnx84;
	wire			Nrnx84;
	wire			Urnx84;
	wire			Bsnx84;
	wire			Isnx84;
	wire			Psnx84;
	wire			Wsnx84;
	wire			Dtnx84;
	wire			Ktnx84;
	wire			Rtnx84;
	wire			Ytnx84;
	wire			Funx84;
	wire			Munx84;
	wire			Tunx84;
	wire			Avnx84;
	wire			Hvnx84;
	wire			Ovnx84;
	wire			Vvnx84;
	wire			Cwnx84;
	wire			Jwnx84;
	wire			Qwnx84;
	wire			Xwnx84;
	wire			Exnx84;
	wire			Lxnx84;
	wire			Sxnx84;
	wire			Zxnx84;
	wire			Gynx84;
	wire			Nynx84;
	wire			Uynx84;
	wire			Bznx84;
	wire			Iznx84;
	wire			Pznx84;
	wire			Wznx84;
	wire			D0ox84;
	wire			K0ox84;
	wire			R0ox84;
	wire			Y0ox84;
	wire			F1ox84;
	wire			M1ox84;
	wire			T1ox84;
	wire			A2ox84;
	wire			H2ox84;
	wire			O2ox84;
	wire			V2ox84;
	wire			C3ox84;
	wire			J3ox84;
	wire			Q3ox84;
	wire			X3ox84;
	wire			E4ox84;
	wire			L4ox84;
	wire			S4ox84;
	wire			Z4ox84;
	wire			G5ox84;
	wire			N5ox84;
	wire			U5ox84;
	wire			B6ox84;
	wire			I6ox84;
	wire			P6ox84;
	wire			W6ox84;
	wire			D7ox84;
	wire			K7ox84;
	wire			R7ox84;
	wire			Y7ox84;
	wire			F8ox84;
	wire			M8ox84;
	wire			T8ox84;
	wire			A9ox84;
	wire			H9ox84;
	wire			O9ox84;
	wire			V9ox84;
	wire			Caox84;
	wire			Jaox84;
	wire			Qaox84;
	wire			Xaox84;
	wire			Ebox84;
	wire			Lbox84;
	wire			Sbox84;
	wire			Zbox84;
	wire			Gcox84;
	wire			Ncox84;
	wire			Ucox84;
	wire			Bdox84;
	wire			Idox84;
	wire			Pdox84;
	wire			Wdox84;
	wire			Deox84;
	wire			Keox84;
	wire			Reox84;
	wire			Yeox84;
	wire			Ffox84;
	wire			Mfox84;
	wire			Tfox84;
	wire			Agox84;
	wire			Hgox84;
	wire			Ogox84;
	wire			Vgox84;
	wire			Chox84;
	wire			Jhox84;
	wire			Qhox84;
	wire			Xhox84;
	wire			Eiox84;
	wire			Liox84;
	wire			Siox84;
	wire			Ziox84;
	wire			Gjox84;
	wire			Njox84;
	wire			Ujox84;
	wire			Bkox84;
	wire			Ikox84;
	wire			Pkox84;
	wire			Wkox84;
	wire			Dlox84;
	wire			Klox84;
	wire			Rlox84;
	wire			Ylox84;
	wire			Fmox84;
	wire			Mmox84;
	wire			Tmox84;
	wire			Anox84;
	wire			Hnox84;
	wire			Onox84;
	wire			Vnox84;
	wire			Coox84;
	wire			Joox84;
	wire			Qoox84;
	wire			Xoox84;
	wire			Epox84;
	wire			Lpox84;
	wire			Spox84;
	wire			Zpox84;
	wire			Gqox84;
	wire			Nqox84;
	wire			Uqox84;
	wire			Brox84;
	wire			Irox84;
	wire			Prox84;
	wire			Wrox84;
	wire			Dsox84;
	wire			Ksox84;
	wire			Rsox84;
	wire			Ysox84;
	wire			Ftox84;
	wire			Mtox84;
	wire			Ttox84;
	wire			Auox84;
	wire			Huox84;
	wire			Ouox84;
	wire			Vuox84;
	wire			Cvox84;
	wire			Jvox84;
	wire			Qvox84;
	wire			Xvox84;
	wire			Ewox84;
	wire			Lwox84;
	wire			Swox84;
	wire			Zwox84;
	wire			Gxox84;
	wire			Nxox84;
	wire			Uxox84;
	wire			Byox84;
	wire			Iyox84;
	wire			Pyox84;
	wire			Wyox84;
	wire			Dzox84;
	wire			Kzox84;
	wire			Rzox84;
	wire			Yzox84;
	wire			F0px84;
	wire			M0px84;
	wire			T0px84;
	wire			A1px84;
	wire			H1px84;
	wire			O1px84;
	wire			V1px84;
	wire			C2px84;
	wire			J2px84;
	wire			Q2px84;
	wire			X2px84;
	wire			E3px84;
	wire			L3px84;
	wire			S3px84;
	wire			Z3px84;
	wire			G4px84;
	wire			N4px84;
	wire			U4px84;
	wire			B5px84;
	wire			I5px84;
	wire			P5px84;
	wire			W5px84;
	wire			D6px84;
	wire			K6px84;
	wire			R6px84;
	wire			Y6px84;
	wire			F7px84;
	wire			M7px84;
	wire			T7px84;
	wire			A8px84;
	wire			H8px84;
	wire			O8px84;
	wire			V8px84;
	wire			C9px84;
	wire			J9px84;
	wire			Q9px84;
	wire			X9px84;
	wire			Eapx84;
	wire			Lapx84;
	wire			Sapx84;
	wire			Zapx84;
	wire			Gbpx84;
	wire			Nbpx84;
	wire			Ubpx84;
	wire			Bcpx84;
	wire			Icpx84;
	wire			Pcpx84;
	wire			Wcpx84;
	wire			Ddpx84;
	wire			Kdpx84;
	wire			Rdpx84;
	wire			Ydpx84;
	wire			Fepx84;
	wire			Mepx84;
	wire			Tepx84;
	wire			Afpx84;
	wire			Hfpx84;
	wire			Ofpx84;
	wire			Vfpx84;
	wire			Cgpx84;
	wire			Jgpx84;
	wire			Qgpx84;
	wire			Xgpx84;
	wire			Ehpx84;
	wire			Lhpx84;
	wire			Shpx84;
	wire			Zhpx84;
	wire			Gipx84;
	wire			Nipx84;
	wire			Uipx84;
	wire			Bjpx84;
	wire			Ijpx84;
	wire			Pjpx84;
	wire			Wjpx84;
	wire			Dkpx84;
	wire			Kkpx84;
	wire			Rkpx84;
	wire			Ykpx84;
	wire			Flpx84;
	wire			Mlpx84;
	wire			Tlpx84;
	wire			Ampx84;
	wire			Hmpx84;
	wire			Ompx84;
	wire			Vmpx84;
	wire			Cnpx84;
	wire			Jnpx84;
	wire			Qnpx84;
	wire			Xnpx84;
	wire			Eopx84;
	wire			Lopx84;
	wire			Sopx84;
	wire			Zopx84;
	wire			Gppx84;
	wire			Nppx84;
	wire			Uppx84;
	wire			Bqpx84;
	wire			Iqpx84;
	wire			Pqpx84;
	wire			Wqpx84;
	wire			Drpx84;
	wire			Krpx84;
	wire			Rrpx84;
	wire			Yrpx84;
	wire			Fspx84;
	wire			Mspx84;
	wire			Tspx84;
	wire			Atpx84;
	wire			Htpx84;
	wire			Otpx84;
	wire			Vtpx84;
	wire			Cupx84;
	wire			Jupx84;
	wire			Qupx84;
	wire			Xupx84;
	wire			Evpx84;
	wire			Lvpx84;
	wire			Svpx84;
	wire			Zvpx84;
	wire			Gwpx84;
	wire			Nwpx84;
	wire			Uwpx84;
	wire			Bxpx84;
	wire			Ixpx84;
	wire			Pxpx84;
	wire			Wxpx84;
	wire			Dypx84;
	wire			Kypx84;
	wire			Rypx84;
	wire			Yypx84;
	wire			Fzpx84;
	wire			Mzpx84;
	wire			Tzpx84;
	wire			A0qx84;
	wire			H0qx84;
	wire			O0qx84;
	wire			V0qx84;
	wire			C1qx84;
	wire			J1qx84;
	wire			Q1qx84;
	wire			X1qx84;
	wire			E2qx84;
	wire			L2qx84;
	wire			S2qx84;
	wire			Z2qx84;
	wire			G3qx84;
	wire			N3qx84;
	wire			U3qx84;
	wire			B4qx84;
	wire			I4qx84;
	wire			P4qx84;
	wire			W4qx84;
	wire			D5qx84;
	wire			K5qx84;
	wire			R5qx84;
	wire			Y5qx84;
	wire			F6qx84;
	wire			M6qx84;
	wire			T6qx84;
	wire			A7qx84;
	wire			H7qx84;
	wire			O7qx84;
	wire			V7qx84;
	wire			C8qx84;
	wire			J8qx84;
	wire			Q8qx84;
	wire			X8qx84;
	wire			E9qx84;
	wire			L9qx84;
	wire			S9qx84;
	wire			Z9qx84;
	wire			Gaqx84;
	wire			Naqx84;
	wire			Uaqx84;
	wire			Bbqx84;
	wire			Ibqx84;
	wire			Pbqx84;
	wire			Wbqx84;
	wire			Dcqx84;
	wire			Kcqx84;
	wire			Rcqx84;
	wire			Ycqx84;
	wire			Fdqx84;
	wire			Mdqx84;
	wire			Tdqx84;
	wire			Aeqx84;
	wire			Heqx84;
	wire			Oeqx84;
	wire			Veqx84;
	wire			Cfqx84;
	wire			Jfqx84;
	wire			Qfqx84;
	wire			Xfqx84;
	wire			Egqx84;
	wire			Lgqx84;
	wire			Sgqx84;
	wire			Zgqx84;
	wire			Ghqx84;
	wire			Nhqx84;
	wire			Uhqx84;
	wire			Biqx84;
	wire			Iiqx84;
	wire			Piqx84;
	wire			Wiqx84;
	wire			Djqx84;
	wire			Kjqx84;
	wire			Rjqx84;
	wire			Yjqx84;
	wire			Fkqx84;
	wire			Mkqx84;
	wire			Tkqx84;
	wire			Alqx84;
	wire			Hlqx84;
	wire			Olqx84;
	wire			Vlqx84;
	wire			Cmqx84;
	wire			Jmqx84;
	wire			Qmqx84;
	wire			Xmqx84;
	wire			Enqx84;
	wire			Lnqx84;
	wire			Snqx84;
	wire			Znqx84;
	wire			Goqx84;
	wire			Noqx84;
	wire			Uoqx84;
	wire			Bpqx84;
	wire			Ipqx84;
	wire			Ppqx84;
	wire			Wpqx84;
	wire			Dqqx84;
	wire			Kqqx84;
	wire			Rqqx84;
	wire			Yqqx84;
	wire			Frqx84;
	wire			Mrqx84;
	wire			Trqx84;
	wire			Asqx84;
	wire			Hsqx84;
	wire			Osqx84;
	wire			Vsqx84;
	wire			Ctqx84;
	wire			Jtqx84;
	wire			Qtqx84;
	wire			Xtqx84;
	wire			Euqx84;
	wire			Luqx84;
	wire			Suqx84;
	wire			Zuqx84;
	wire			Gvqx84;
	wire			Nvqx84;
	wire			Uvqx84;
	wire			Bwqx84;
	wire			Iwqx84;
	wire			Pwqx84;
	wire			Wwqx84;
	wire			Dxqx84;
	wire			Kxqx84;
	wire			Rxqx84;
	wire			Yxqx84;
	wire			Fyqx84;
	wire			Myqx84;
	wire			Tyqx84;
	wire			Azqx84;
	wire			Hzqx84;
	wire			Ozqx84;
	wire			Vzqx84;
	wire			C0rx84;
	wire			J0rx84;
	wire			Q0rx84;
	wire			X0rx84;
	wire			E1rx84;
	wire			L1rx84;
	wire			S1rx84;
	wire			Z1rx84;
	wire			G2rx84;
	wire			N2rx84;
	wire			U2rx84;
	wire			B3rx84;
	wire			I3rx84;
	wire			P3rx84;
	wire			W3rx84;
	wire			D4rx84;
	wire			K4rx84;
	wire			R4rx84;
	wire			Y4rx84;
	wire			F5rx84;
	wire			M5rx84;
	wire			T5rx84;
	wire			A6rx84;
	wire			H6rx84;
	wire			O6rx84;
	wire			V6rx84;
	wire			C7rx84;
	wire			J7rx84;
	wire			Q7rx84;
	wire			X7rx84;
	wire			E8rx84;
	wire			L8rx84;
	wire			S8rx84;
	wire			Z8rx84;
	wire			G9rx84;
	wire			N9rx84;
	wire			U9rx84;
	wire			Barx84;
	wire			Iarx84;
	wire			Parx84;
	wire			Warx84;
	wire			Dbrx84;
	wire			Kbrx84;
	wire			Rbrx84;
	wire			Ybrx84;
	wire			Fcrx84;
	wire			Mcrx84;
	wire			Tcrx84;
	wire			Adrx84;
	wire			Hdrx84;
	wire			Odrx84;
	wire			Vdrx84;
	wire			Cerx84;
	wire			Jerx84;
	wire			Qerx84;
	wire			Xerx84;
	wire			Efrx84;
	wire			Lfrx84;
	wire			Sfrx84;
	wire			Zfrx84;
	wire			Ggrx84;
	wire			Ngrx84;
	wire			Ugrx84;
	wire			Bhrx84;
	wire			Ihrx84;
	wire			Phrx84;
	wire			Whrx84;
	wire			Dirx84;
	wire			Kirx84;
	wire			Rirx84;
	wire			Yirx84;
	wire			Fjrx84;
	wire			Mjrx84;
	wire			Tjrx84;
	wire			Akrx84;
	wire			Hkrx84;
	wire			Okrx84;
	wire			Vkrx84;
	wire			Clrx84;
	wire			Jlrx84;
	wire			Qlrx84;
	wire			Xlrx84;
	wire			Emrx84;
	wire			Lmrx84;
	wire			Smrx84;
	wire			Zmrx84;
	wire			Gnrx84;
	wire			Nnrx84;
	wire			Unrx84;
	wire			Borx84;
	wire			Iorx84;
	wire			Porx84;
	wire			Worx84;
	wire			Dprx84;
	wire			Kprx84;
	wire			Rprx84;
	wire			Yprx84;
	wire			Fqrx84;
	wire			Mqrx84;
	wire			Tqrx84;
	wire			Arrx84;
	wire			Hrrx84;
	wire			Orrx84;
	wire			Vrrx84;
	wire			Csrx84;
	wire			Jsrx84;
	wire			Qsrx84;
	wire			Xsrx84;
	wire			Etrx84;
	wire			Ltrx84;
	wire			Strx84;
	wire			Ztrx84;
	wire			Gurx84;
	wire			Nurx84;
	wire			Uurx84;
	wire			Bvrx84;
	wire			Ivrx84;
	wire			Pvrx84;
	wire			Wvrx84;
	wire			Dwrx84;
	wire			Kwrx84;
	wire			Rwrx84;
	wire			Ywrx84;
	wire			Fxrx84;
	wire			Mxrx84;
	wire			Txrx84;
	wire			Ayrx84;
	wire			Hyrx84;
	wire			Oyrx84;
	wire			Vyrx84;
	wire			Czrx84;
	wire			Jzrx84;
	wire			Qzrx84;
	wire			Xzrx84;
	wire			E0sx84;
	wire			L0sx84;
	wire			S0sx84;
	wire			Z0sx84;
	wire			G1sx84;
	wire			N1sx84;
	wire			U1sx84;
	wire			B2sx84;
	wire			I2sx84;
	wire			P2sx84;
	wire			W2sx84;
	wire			D3sx84;
	wire			K3sx84;
	wire			R3sx84;
	wire			Y3sx84;
	wire			F4sx84;
	wire			M4sx84;
	wire			T4sx84;
	wire			A5sx84;
	wire			H5sx84;
	wire			O5sx84;
	wire			V5sx84;
	wire			C6sx84;
	wire			J6sx84;
	wire			Q6sx84;
	wire			X6sx84;
	wire			E7sx84;
	wire			L7sx84;
	wire			S7sx84;
	wire			Z7sx84;
	wire			G8sx84;
	wire			N8sx84;
	wire			U8sx84;
	wire			B9sx84;
	wire			I9sx84;
	wire			P9sx84;
	wire			W9sx84;
	wire			Dasx84;
	wire			Kasx84;
	wire			Rasx84;
	wire			Yasx84;
	wire			Fbsx84;
	wire			Mbsx84;
	wire			Tbsx84;
	wire			Acsx84;
	wire			Hcsx84;
	wire			Ocsx84;
	wire			Vcsx84;
	wire			Cdsx84;
	wire			Jdsx84;
	wire			Qdsx84;
	wire			Xdsx84;
	wire			Eesx84;
	wire			Lesx84;
	wire			Sesx84;
	wire			Zesx84;
	wire			Gfsx84;
	wire			Nfsx84;
	wire			Ufsx84;
	wire			Bgsx84;
	wire			Igsx84;
	wire			Pgsx84;
	wire			Wgsx84;
	wire			Dhsx84;
	wire			Khsx84;
	wire			Rhsx84;
	wire			Yhsx84;
	wire			Fisx84;
	wire			Misx84;
	wire			Tisx84;
	wire			Ajsx84;
	wire			Hjsx84;
	wire			Ojsx84;
	wire			Vjsx84;
	wire			Cksx84;
	wire			Jksx84;
	wire			Qksx84;
	wire			Xksx84;
	wire			Elsx84;
	wire			Llsx84;
	wire			Slsx84;
	wire			Zlsx84;
	wire			Gmsx84;
	wire			Nmsx84;
	wire			Umsx84;
	wire			Bnsx84;
	wire			Insx84;
	wire			Pnsx84;
	wire			Wnsx84;
	wire			Dosx84;
	wire			Kosx84;
	wire			Rosx84;
	wire			Yosx84;
	wire			Fpsx84;
	wire			Mpsx84;
	wire			Tpsx84;
	wire			Aqsx84;
	wire			Hqsx84;
	wire			Oqsx84;
	wire			Vqsx84;
	wire			Crsx84;
	wire			Jrsx84;
	wire			Qrsx84;
	wire			Xrsx84;
	wire			Essx84;
	wire			Lssx84;
	wire			Sssx84;
	wire			Zssx84;
	wire			Gtsx84;
	wire			Ntsx84;
	wire			Utsx84;
	wire			Busx84;
	wire			Iusx84;
	wire			Pusx84;
	wire			Wusx84;
	wire			Dvsx84;
	wire			Kvsx84;
	wire			Rvsx84;
	wire			Yvsx84;
	wire			Fwsx84;
	wire			Mwsx84;
	wire			Twsx84;
	wire			Axsx84;
	wire			Hxsx84;
	wire			Oxsx84;
	wire			Vxsx84;
	wire			Cysx84;
	wire			Jysx84;
	wire			Qysx84;
	wire			Xysx84;
	wire			Ezsx84;
	wire			Lzsx84;
	wire			Szsx84;
	wire			Zzsx84;
	wire			G0tx84;
	wire			N0tx84;
	wire			U0tx84;
	wire			B1tx84;
	wire			I1tx84;
	wire			P1tx84;
	wire			W1tx84;
	wire			D2tx84;
	wire			K2tx84;
	wire			R2tx84;
	wire			Y2tx84;
	wire			F3tx84;
	wire			M3tx84;
	wire			T3tx84;
	wire			A4tx84;
	wire			H4tx84;
	wire			O4tx84;
	wire			V4tx84;
	wire			C5tx84;
	wire			J5tx84;
	wire			Q5tx84;
	wire			X5tx84;
	wire			E6tx84;
	wire			L6tx84;
	wire			S6tx84;
	wire			Z6tx84;
	wire			G7tx84;
	wire			N7tx84;
	wire			U7tx84;
	wire			B8tx84;
	wire			I8tx84;
	wire			P8tx84;
	wire			W8tx84;
	wire			D9tx84;
	wire			K9tx84;
	wire			R9tx84;
	wire			Y9tx84;
	wire			Fatx84;
	wire			Matx84;
	wire			Tatx84;
	wire			Abtx84;
	wire			Hbtx84;
	wire			Obtx84;
	wire			Vbtx84;
	wire			Cctx84;
	wire			Jctx84;
	wire			Qctx84;
	wire			Xctx84;
	wire			Edtx84;
	wire			Ldtx84;
	wire			Sdtx84;
	wire			Zdtx84;
	wire			Getx84;
	wire			Netx84;
	wire			Uetx84;
	wire			Bftx84;
	wire			Iftx84;
	wire			Pftx84;
	wire			Wftx84;
	wire			Dgtx84;
	wire			Kgtx84;
	wire			Rgtx84;
	wire			Ygtx84;
	wire			Fhtx84;
	wire			Mhtx84;
	wire			Thtx84;
	wire			Aitx84;
	wire			Hitx84;
	wire			Oitx84;
	wire			Vitx84;
	wire			Cjtx84;
	wire			Jjtx84;
	wire			Qjtx84;
	wire			Xjtx84;
	wire			Ektx84;
	wire			Lktx84;
	wire			Sktx84;
	wire			Zktx84;
	wire			Gltx84;
	wire			Nltx84;
	wire			Ultx84;
	wire			Bmtx84;
	wire			Imtx84;
	wire			Pmtx84;
	wire			Wmtx84;
	wire			Dntx84;
	wire			Kntx84;
	wire			Rntx84;
	wire			Yntx84;
	wire			Fotx84;
	wire			Motx84;
	wire			Totx84;
	wire			Aptx84;
	wire			Hptx84;
	wire			Optx84;
	wire			Vptx84;
	wire			Cqtx84;
	wire			Jqtx84;
	wire			Qqtx84;
	wire			Xqtx84;
	wire			Ertx84;
	wire			Lrtx84;
	wire			Srtx84;
	wire			Zrtx84;
	wire			Gstx84;
	wire			Nstx84;
	wire			Ustx84;
	wire			Bttx84;
	wire			Ittx84;
	wire			Pttx84;
	wire			Wttx84;
	wire			Dutx84;
	wire			Kutx84;
	wire			Rutx84;
	wire			Yutx84;
	wire			Fvtx84;
	wire			Mvtx84;
	wire			Tvtx84;
	wire			Awtx84;
	wire			Hwtx84;
	wire			Owtx84;
	wire			Vwtx84;
	wire			Cxtx84;
	wire			Jxtx84;
	wire			Qxtx84;
	wire			Xxtx84;
	wire			Eytx84;
	wire			Lytx84;
	wire			Sytx84;
	wire			Zytx84;
	wire			Gztx84;
	wire			Nztx84;
	wire			Uztx84;
	wire			B0ux84;
	wire			I0ux84;
	wire			P0ux84;
	wire			W0ux84;
	wire			D1ux84;
	wire			K1ux84;
	wire			R1ux84;
	wire			Y1ux84;
	wire			F2ux84;
	wire			M2ux84;
	wire			T2ux84;
	wire			A3ux84;
	wire			H3ux84;
	wire			O3ux84;
	wire			V3ux84;
	wire			C4ux84;
	wire			J4ux84;
	wire			Q4ux84;
	wire			X4ux84;
	wire			E5ux84;
	wire			L5ux84;
	wire			S5ux84;
	wire			Z5ux84;
	wire			G6ux84;
	wire			N6ux84;
	wire			U6ux84;
	wire			B7ux84;
	wire			I7ux84;
	wire			P7ux84;
	wire			W7ux84;
	wire			D8ux84;
	wire			K8ux84;
	wire			R8ux84;
	wire			Y8ux84;
	wire			F9ux84;
	wire			M9ux84;
	wire			T9ux84;
	wire			Aaux84;
	wire			Haux84;
	wire			Oaux84;
	wire			Vaux84;
	wire			Cbux84;
	wire			Jbux84;
	wire			Qbux84;
	wire			Xbux84;
	wire			Ecux84;
	wire			Lcux84;
	wire			Scux84;
	wire			Zcux84;
	wire			Gdux84;
	wire			Ndux84;
	wire			Udux84;
	wire			Beux84;
	wire			Ieux84;
	wire			Peux84;
	wire			Weux84;
	wire			Dfux84;
	wire			Kfux84;
	wire			Rfux84;
	wire			Yfux84;
	wire			Fgux84;
	wire			Mgux84;
	wire			Tgux84;
	wire			Ahux84;
	wire			Hhux84;
	wire			Ohux84;
	wire			Vhux84;
	wire			Ciux84;
	wire			Jiux84;
	wire			Qiux84;
	wire			Xiux84;
	wire			Ejux84;
	wire			Ljux84;
	wire			Sjux84;
	wire			Zjux84;
	wire			Gkux84;
	wire			Nkux84;
	wire			Ukux84;
	wire			Blux84;
	wire			Ilux84;
	wire			Plux84;
	wire			Wlux84;
	wire			Dmux84;
	wire			Kmux84;
	wire			Rmux84;
	wire			Ymux84;
	wire			Fnux84;
	wire			Mnux84;
	wire			Tnux84;
	wire			Aoux84;
	wire			Houx84;
	wire			Ooux84;
	wire			Voux84;
	wire			Cpux84;
	wire			Jpux84;
	wire			Qpux84;
	wire			Xpux84;
	wire			Equx84;
	wire			Lqux84;
	wire			Squx84;
	wire			Zqux84;
	wire			Grux84;
	wire			Nrux84;
	wire			Urux84;
	wire			Bsux84;
	wire			Isux84;
	wire			Psux84;
	wire			Wsux84;
	wire			Dtux84;
	wire			Ktux84;
	wire			Rtux84;
	wire			Ytux84;
	wire			Fuux84;
	wire			Muux84;
	wire			Tuux84;
	wire			Avux84;
	wire			Hvux84;
	wire			Ovux84;
	wire			Vvux84;
	wire			Cwux84;
	wire			Jwux84;
	wire			Qwux84;
	wire			Xwux84;
	wire			Exux84;
	wire			Lxux84;
	wire			Sxux84;
	wire			Zxux84;
	wire			Gyux84;
	wire			Nyux84;
	wire			Uyux84;
	wire			Bzux84;
	wire			Izux84;
	wire			Pzux84;
	wire			Wzux84;
	wire			D0vx84;
	wire			K0vx84;
	wire			R0vx84;
	wire			Y0vx84;
	wire			F1vx84;
	wire			M1vx84;
	wire			T1vx84;
	wire			A2vx84;
	wire			H2vx84;
	wire			O2vx84;
	wire			V2vx84;
	wire			C3vx84;
	wire			J3vx84;
	wire			Q3vx84;
	wire			X3vx84;
	wire			E4vx84;
	wire			L4vx84;
	wire			S4vx84;
	wire			Z4vx84;
	wire			G5vx84;
	wire			N5vx84;
	wire			U5vx84;
	wire			B6vx84;
	wire			I6vx84;
	wire			P6vx84;
	wire			W6vx84;
	wire			D7vx84;
	wire			K7vx84;
	wire			R7vx84;
	wire			Y7vx84;
	wire			F8vx84;
	wire			M8vx84;
	wire			T8vx84;
	wire			A9vx84;
	wire			H9vx84;
	wire			O9vx84;
	wire			V9vx84;
	wire			Cavx84;
	wire			Javx84;
	wire			Qavx84;
	wire			Xavx84;
	wire			Ebvx84;
	wire			Lbvx84;
	wire			Sbvx84;
	wire			Zbvx84;
	wire			Gcvx84;
	wire			Ncvx84;
	wire			Ucvx84;
	wire			Bdvx84;
	wire			Idvx84;
	wire			Pdvx84;
	wire			Wdvx84;
	wire			Devx84;
	wire			Kevx84;
	wire			Revx84;
	wire			Yevx84;
	wire			Ffvx84;
	wire			Mfvx84;
	wire			Tfvx84;
	wire			Agvx84;
	wire			Hgvx84;
	wire			Ogvx84;
	wire			Vgvx84;
	wire			Chvx84;
	wire			Jhvx84;
	wire			Qhvx84;
	wire			Xhvx84;
	wire			Eivx84;
	wire			Livx84;
	wire			Sivx84;
	wire			Zivx84;
	wire			Gjvx84;
	wire			Njvx84;
	wire			Ujvx84;
	wire			Bkvx84;
	wire			Ikvx84;
	wire			Pkvx84;
	wire			Wkvx84;
	wire			Dlvx84;
	wire			Klvx84;
	wire			Rlvx84;
	wire			Ylvx84;
	wire			Fmvx84;
	wire			Mmvx84;
	wire			Tmvx84;
	wire			Anvx84;
	wire			Hnvx84;
	wire			Onvx84;
	wire			Vnvx84;
	wire			Covx84;
	wire			Jovx84;
	wire			Qovx84;
	wire			Xovx84;
	wire			Epvx84;
	wire			Lpvx84;
	wire			Spvx84;
	wire			Zpvx84;
	wire			Gqvx84;
	wire			Nqvx84;
	wire			Uqvx84;
	wire			Brvx84;
	wire			Irvx84;
	wire			Prvx84;
	wire			Wrvx84;
	wire			Dsvx84;
	wire			Ksvx84;
	wire			Rsvx84;
	wire			Ysvx84;
	wire			Ftvx84;
	wire			Mtvx84;
	wire			Ttvx84;
	wire			Auvx84;
	wire			Huvx84;
	wire			Ouvx84;
	wire			Vuvx84;
	wire			Cvvx84;
	wire			Jvvx84;
	wire			Qvvx84;
	wire			Xvvx84;
	wire			Ewvx84;
	wire			Lwvx84;
	wire			Swvx84;
	wire			Zwvx84;
	wire			Gxvx84;
	wire			Nxvx84;
	wire			Uxvx84;
	wire			Byvx84;
	wire			Iyvx84;
	wire			Pyvx84;
	wire			Wyvx84;
	wire			Dzvx84;
	wire			Kzvx84;
	wire			Rzvx84;
	wire			Yzvx84;
	wire			F0wx84;
	wire			M0wx84;
	wire			T0wx84;
	wire			A1wx84;
	wire			H1wx84;
	wire			O1wx84;
	wire			V1wx84;
	wire			C2wx84;
	wire			J2wx84;
	wire			Q2wx84;
	wire			X2wx84;
	wire			E3wx84;
	wire			L3wx84;
	wire			S3wx84;
	wire			Z3wx84;
	wire			G4wx84;
	wire			N4wx84;
	wire			U4wx84;
	wire			B5wx84;
	wire			I5wx84;
	wire			P5wx84;
	wire			W5wx84;
	wire			D6wx84;
	wire			K6wx84;
	wire			R6wx84;
	wire			Y6wx84;
	wire			F7wx84;
	wire			M7wx84;
	wire			T7wx84;
	wire			A8wx84;
	wire			H8wx84;
	wire			O8wx84;
	wire			V8wx84;
	wire			C9wx84;
	wire			J9wx84;
	wire			Q9wx84;
	wire			X9wx84;
	wire			Eawx84;
	wire			Lawx84;
	wire			Sawx84;
	wire			Zawx84;
	wire			Gbwx84;
	wire			Nbwx84;
	wire			Ubwx84;
	wire			Bcwx84;
	wire			Icwx84;
	wire			Pcwx84;
	wire			Wcwx84;
	wire			Ddwx84;
	wire			Kdwx84;
	wire			Rdwx84;
	wire			Ydwx84;
	wire			Fewx84;
	wire			Mewx84;
	wire			Tewx84;
	wire			Afwx84;
	wire			Hfwx84;
	wire			Ofwx84;
	wire			Vfwx84;
	wire			Cgwx84;
	wire			Jgwx84;
	wire			Qgwx84;
	wire			Xgwx84;
	wire			Ehwx84;
	wire			Lhwx84;
	wire			Shwx84;
	wire			Zhwx84;
	wire			Giwx84;
	wire			Niwx84;
	wire			Uiwx84;
	wire			Bjwx84;
	wire			Ijwx84;
	wire			Pjwx84;
	wire			Wjwx84;
	wire			Dkwx84;
	wire			Kkwx84;
	wire			Rkwx84;
	wire			Ykwx84;
	wire			Flwx84;
	wire			Mlwx84;
	wire			Tlwx84;
	wire			Amwx84;
	wire			Hmwx84;
	wire			Omwx84;
	wire			Vmwx84;
	wire			Cnwx84;
	wire			Jnwx84;
	wire			Qnwx84;
	wire			Xnwx84;
	wire			Eowx84;
	wire			Lowx84;
	wire			Sowx84;
	wire			Zowx84;
	wire			Gpwx84;
	wire			Npwx84;
	wire			Upwx84;
	wire			Bqwx84;
	wire			Iqwx84;
	wire			Pqwx84;
	wire			Wqwx84;
	wire			Drwx84;
	wire			Krwx84;
	wire			Rrwx84;
	wire			Yrwx84;
	wire			Fswx84;
	wire			Mswx84;
	wire			Tswx84;
	wire			Atwx84;
	wire			Htwx84;
	wire			Otwx84;
	wire			Vtwx84;
	wire			Cuwx84;
	wire			Juwx84;
	wire			Quwx84;
	wire			Xuwx84;
	wire			Evwx84;
	wire			Lvwx84;
	wire			Svwx84;
	wire			Zvwx84;
	wire			Gwwx84;
	wire			Nwwx84;
	wire			Uwwx84;
	wire			Bxwx84;
	wire			Ixwx84;
	wire			Pxwx84;
	wire			Wxwx84;
	wire			Dywx84;
	wire			Kywx84;
	wire			Rywx84;
	wire			Yywx84;
	wire			Fzwx84;
	wire			Mzwx84;
	wire			Tzwx84;
	wire			A0xx84;
	wire			H0xx84;
	wire			O0xx84;
	wire			V0xx84;
	wire			C1xx84;
	wire			J1xx84;
	wire			Q1xx84;
	wire			X1xx84;
	wire			E2xx84;
	wire			L2xx84;
	wire			S2xx84;
	wire			Z2xx84;
	wire			G3xx84;
	wire			N3xx84;
	wire			U3xx84;
	wire			B4xx84;
	wire			I4xx84;
	wire			P4xx84;
	wire			W4xx84;
	wire			D5xx84;
	wire			K5xx84;
	wire			R5xx84;
	wire			Y5xx84;
	wire			F6xx84;
	wire			M6xx84;
	wire			T6xx84;
	wire			A7xx84;
	wire			H7xx84;
	wire			O7xx84;
	wire			V7xx84;
	wire			C8xx84;
	wire			J8xx84;
	wire			Q8xx84;
	wire			X8xx84;
	wire			E9xx84;
	wire			L9xx84;
	wire			S9xx84;
	wire			Z9xx84;
	wire			Gaxx84;
	wire			Naxx84;
	wire			Uaxx84;
	wire			Bbxx84;
	wire			Ibxx84;
	wire			Pbxx84;
	wire			Wbxx84;
	wire			Dcxx84;
	wire			Kcxx84;
	wire			Rcxx84;
	wire			Ycxx84;
	wire			Fdxx84;
	wire			Mdxx84;
	wire			Tdxx84;
	wire			Aexx84;
	wire			Hexx84;
	wire			Oexx84;
	wire			Vexx84;
	wire			Cfxx84;
	wire			Jfxx84;
	wire			Qfxx84;
	wire			Xfxx84;
	wire			Egxx84;
	wire			Lgxx84;
	wire			Sgxx84;
	wire			Zgxx84;
	wire			Ghxx84;
	wire			Nhxx84;
	wire			Uhxx84;
	wire			Bixx84;
	wire			Iixx84;
	wire			Pixx84;
	wire			Wixx84;
	wire			Djxx84;
	wire			Kjxx84;
	wire			Rjxx84;
	wire			Yjxx84;
	wire			Fkxx84;
	wire			Mkxx84;
	wire			Tkxx84;
	wire			Alxx84;
	wire			Hlxx84;
	wire			Olxx84;
	wire			Vlxx84;
	wire			Cmxx84;
	wire			Jmxx84;
	wire			Qmxx84;
	wire			Xmxx84;
	wire			Enxx84;
	wire			Lnxx84;
	wire			Snxx84;
	wire			Znxx84;
	wire			Goxx84;
	wire			Noxx84;
	wire			Uoxx84;
	wire			Bpxx84;
	wire			Ipxx84;
	wire			Ppxx84;
	wire			Wpxx84;
	wire			Dqxx84;
	wire			Kqxx84;
	wire			Rqxx84;
	wire			Yqxx84;
	wire			Frxx84;
	wire			Mrxx84;
	wire			Trxx84;
	wire			Asxx84;
	wire			Hsxx84;
	wire			Osxx84;
	wire			Vsxx84;
	wire			Ctxx84;
	wire			Jtxx84;
	wire			Qtxx84;
	wire			Xtxx84;
	wire			Euxx84;
	wire			Luxx84;
	wire			Suxx84;
	wire			Zuxx84;
	wire			Gvxx84;
	wire			Nvxx84;
	wire			Uvxx84;
	wire			Bwxx84;
	wire			Iwxx84;
	wire			Pwxx84;
	wire			Wwxx84;
	wire			Dxxx84;
	wire			Kxxx84;
	wire			Rxxx84;
	wire			Yxxx84;
	wire			Fyxx84;
	wire			Myxx84;
	wire			Tyxx84;
	wire			Azxx84;
	wire			Hzxx84;
	wire			Ozxx84;
	wire			Vzxx84;
	wire			C0yx84;
	wire			J0yx84;
	wire			Q0yx84;
	wire			X0yx84;
	wire			E1yx84;
	wire			L1yx84;
	wire			S1yx84;
	wire			Z1yx84;
	wire			G2yx84;
	wire			N2yx84;
	wire			U2yx84;
	wire			B3yx84;
	wire			I3yx84;
	wire			P3yx84;
	wire			W3yx84;
	wire			D4yx84;
	wire			K4yx84;
	wire			R4yx84;
	wire			Y4yx84;
	wire			F5yx84;
	wire			M5yx84;
	wire			T5yx84;
	wire			A6yx84;
	wire			H6yx84;
	wire			O6yx84;
	wire			V6yx84;
	wire			C7yx84;
	wire			J7yx84;
	wire			Q7yx84;
	wire			X7yx84;
	wire			E8yx84;
	wire			L8yx84;
	wire			S8yx84;
	wire			Z8yx84;
	wire			G9yx84;
	wire			N9yx84;
	wire			U9yx84;
	wire			Bayx84;
	wire			Iayx84;
	wire			Payx84;
	wire			Wayx84;
	wire			Dbyx84;
	wire			Kbyx84;
	wire			Rbyx84;
	wire			Ybyx84;
	wire			Fcyx84;
	wire			Mcyx84;
	wire			Tcyx84;
	wire			Adyx84;
	wire			Hdyx84;
	wire			Odyx84;
	wire			Vdyx84;
	wire			Ceyx84;
	wire			Jeyx84;
	wire			Qeyx84;
	wire			Xeyx84;
	wire			Efyx84;
	wire			Lfyx84;
	wire			Sfyx84;
	wire			Zfyx84;
	wire			Ggyx84;
	wire			Ngyx84;
	wire			Ugyx84;
	wire			Bhyx84;
	wire			Ihyx84;
	wire			Phyx84;
	wire			Whyx84;
	wire			Diyx84;
	wire			Kiyx84;
	wire			Riyx84;
	wire			Yiyx84;
	wire			Fjyx84;
	wire			Mjyx84;
	wire			Tjyx84;
	wire			Akyx84;
	wire			Hkyx84;
	wire			Okyx84;
	wire			Vkyx84;
	wire			Clyx84;
	wire			Jlyx84;
	wire			Qlyx84;
	wire			Xlyx84;
	wire			Emyx84;
	wire			Lmyx84;
	wire			Smyx84;
	wire			Zmyx84;
	wire			Gnyx84;
	wire			Nnyx84;
	wire			Unyx84;
	wire			Boyx84;
	wire			Ioyx84;
	wire			Poyx84;
	wire			Woyx84;
	wire			Dpyx84;
	wire			Kpyx84;
	wire			Rpyx84;
	wire			Ypyx84;
	wire			Fqyx84;
	wire			Mqyx84;
	wire			Tqyx84;
	wire			Aryx84;
	wire			Hryx84;
	wire			Oryx84;
	wire			Vryx84;
	wire			Csyx84;
	wire			Jsyx84;
	wire			Qsyx84;
	wire			Xsyx84;
	wire			Etyx84;
	wire			Ltyx84;
	wire			Styx84;
	wire			Ztyx84;
	wire			Guyx84;
	wire			Nuyx84;
	wire			Uuyx84;
	wire			Bvyx84;
	wire			Ivyx84;
	wire			Pvyx84;
	wire			Wvyx84;
	wire			Dwyx84;
	wire			Kwyx84;
	wire			Rwyx84;
	wire			Ywyx84;
	wire			Fxyx84;
	wire			Mxyx84;
	wire			Txyx84;
	wire			Ayyx84;
	wire			Hyyx84;
	wire			Oyyx84;
	wire			Vyyx84;
	wire			Czyx84;
	wire			Jzyx84;
	wire			Qzyx84;
	wire			Xzyx84;
	wire			E0zx84;
	wire			L0zx84;
	wire			S0zx84;
	wire			Z0zx84;
	wire			G1zx84;
	wire			N1zx84;
	wire			U1zx84;
	wire			B2zx84;
	wire			I2zx84;
	wire			P2zx84;
	wire			W2zx84;
	wire			D3zx84;
	wire			K3zx84;
	wire			R3zx84;
	wire			Y3zx84;
	wire			F4zx84;
	wire			M4zx84;
	wire			T4zx84;
	wire			A5zx84;
	wire			H5zx84;
	wire			O5zx84;
	wire			V5zx84;
	wire			C6zx84;
	wire			J6zx84;
	wire			Q6zx84;
	wire			X6zx84;
	wire			E7zx84;
	wire			L7zx84;
	wire			S7zx84;
	wire			Z7zx84;
	wire			G8zx84;
	wire			N8zx84;
	wire			U8zx84;
	wire			B9zx84;
	wire			I9zx84;
	wire			P9zx84;
	wire			W9zx84;
	wire			Dazx84;
	wire			Kazx84;
	wire			Razx84;
	wire			Yazx84;
	wire			Fbzx84;
	wire			Mbzx84;
	wire			Tbzx84;
	wire			Aczx84;
	wire			Hczx84;
	wire			Oczx84;
	wire			Vczx84;
	wire			Cdzx84;
	wire			Jdzx84;
	wire			Qdzx84;
	wire			Xdzx84;
	wire			Eezx84;
	wire			Lezx84;
	wire			Sezx84;
	wire			Zezx84;
	wire			Gfzx84;
	wire			Nfzx84;
	wire			Ufzx84;
	wire			Bgzx84;
	wire			Igzx84;
	wire			Pgzx84;
	wire			Wgzx84;
	wire			Dhzx84;
	wire			Khzx84;
	wire			Rhzx84;
	wire			Yhzx84;
	wire			Fizx84;
	wire			Mizx84;
	wire			Tizx84;
	wire			Ajzx84;
	wire			Hjzx84;
	wire			Ojzx84;
	wire			Vjzx84;
	wire			Ckzx84;
	wire			Jkzx84;
	wire			Qkzx84;
	wire			Xkzx84;
	wire			Elzx84;
	wire			Llzx84;
	wire			Slzx84;
	wire			Zlzx84;
	wire			Gmzx84;
	wire			Nmzx84;
	wire			Umzx84;
	wire			Bnzx84;
	wire			Inzx84;
	wire			Pnzx84;
	wire			Wnzx84;
	wire			Dozx84;
	wire			Kozx84;
	wire			Rozx84;
	wire			Yozx84;
	wire			Fpzx84;
	wire			Mpzx84;
	wire			Tpzx84;
	wire			Aqzx84;
	wire			Hqzx84;
	wire			Oqzx84;
	wire			Vqzx84;
	wire			Crzx84;
	wire			Jrzx84;
	wire			Qrzx84;
	wire			Xrzx84;
	wire			Eszx84;
	wire			Lszx84;
	wire			Sszx84;
	wire			Zszx84;
	wire			Gtzx84;
	wire			Ntzx84;
	wire			Utzx84;
	wire			Buzx84;
	wire			Iuzx84;
	wire			Puzx84;
	wire			Wuzx84;
	wire			Dvzx84;
	wire			Kvzx84;
	wire			Rvzx84;
	wire			Yvzx84;
	wire			Fwzx84;
	wire			Mwzx84;
	wire			Twzx84;
	wire			Axzx84;
	wire			Hxzx84;
	wire			Oxzx84;
	wire			Vxzx84;
	wire			Cyzx84;
	wire			Jyzx84;
	wire			Qyzx84;
	wire			Xyzx84;
	wire			Ezzx84;
	wire			Lzzx84;
	wire			Szzx84;
	wire			Zzzx84;
	wire			G00y84;
	wire			N00y84;
	wire			U00y84;
	wire			B10y84;
	wire			I10y84;
	wire			P10y84;
	wire			W10y84;
	wire			D20y84;
	wire			K20y84;
	wire			R20y84;
	wire			Y20y84;
	wire			F30y84;
	wire			M30y84;
	wire			T30y84;
	wire			A40y84;
	wire			H40y84;
	wire			O40y84;
	wire			V40y84;
	wire			C50y84;
	wire			J50y84;
	wire			Q50y84;
	wire			X50y84;
	wire			E60y84;
	wire			L60y84;
	wire			S60y84;
	wire			Z60y84;
	wire			G70y84;
	wire			N70y84;
	wire			U70y84;
	wire			B80y84;
	wire			I80y84;
	wire			P80y84;
	wire			W80y84;
	wire			D90y84;
	wire			K90y84;
	wire			R90y84;
	wire			Y90y84;
	wire			Fa0y84;
	wire			Ma0y84;
	wire			Ta0y84;
	wire			Ab0y84;
	wire			Hb0y84;
	wire			Ob0y84;
	wire			Vb0y84;
	wire			Cc0y84;
	wire			Jc0y84;
	wire			Qc0y84;
	wire			Xc0y84;
	wire			Ed0y84;
	wire			Ld0y84;
	wire			Sd0y84;
	wire			Zd0y84;
	wire			Ge0y84;
	wire			Ne0y84;
	wire			Ue0y84;
	wire			Bf0y84;
	wire			If0y84;
	wire			Pf0y84;
	wire			Wf0y84;
	wire			Dg0y84;
	wire			Kg0y84;
	wire			Rg0y84;
	wire			Yg0y84;
	wire			Fh0y84;
	wire			Mh0y84;
	wire			Th0y84;
	wire			Ai0y84;
	wire			Hi0y84;
	wire			Oi0y84;
	wire			Vi0y84;
	wire			Cj0y84;
	wire			Jj0y84;
	wire			Qj0y84;
	wire			Xj0y84;
	wire			Ek0y84;
	wire			Lk0y84;
	wire			Sk0y84;
	wire			Zk0y84;
	wire			Gl0y84;
	wire			Nl0y84;
	wire			Ul0y84;
	wire			Bm0y84;
	wire			Im0y84;
	wire			Pm0y84;
	wire			Wm0y84;
	wire			Dn0y84;
	wire			Kn0y84;
	wire			Rn0y84;
	wire			Yn0y84;
	wire			Fo0y84;
	wire			Mo0y84;
	wire			To0y84;
	wire			Ap0y84;
	wire			Hp0y84;
	wire			Op0y84;
	wire			Vp0y84;
	wire			Cq0y84;
	wire			Jq0y84;
	wire			Qq0y84;
	wire			Xq0y84;
	wire			Er0y84;
	wire			Lr0y84;
	wire			Sr0y84;
	wire			Zr0y84;
	wire			Gs0y84;
	wire			Ns0y84;
	wire			Us0y84;
	wire			Bt0y84;
	wire			It0y84;
	wire			Pt0y84;
	wire			Wt0y84;
	wire			Du0y84;
	wire			Ku0y84;
	wire			Ru0y84;
	wire			Yu0y84;
	wire			Fv0y84;
	wire			Mv0y84;
	wire			Tv0y84;
	wire			Aw0y84;
	wire			Hw0y84;
	wire			Ow0y84;
	wire			Vw0y84;
	wire			Cx0y84;
	wire			Jx0y84;
	wire			Qx0y84;
	wire			Xx0y84;
	wire			Ey0y84;
	wire			Ly0y84;
	wire			Sy0y84;
	wire			Zy0y84;
	wire			Gz0y84;
	wire			Nz0y84;
	wire			Uz0y84;
	wire			B01y84;
	wire			I01y84;
	wire			P01y84;
	wire			W01y84;
	wire			D11y84;
	wire			K11y84;
	wire			R11y84;
	wire			Y11y84;
	wire			F21y84;
	wire			M21y84;
	wire			T21y84;
	wire			A31y84;
	wire			H31y84;
	wire			O31y84;
	wire			V31y84;
	wire			C41y84;
	wire			J41y84;
	wire			Q41y84;
	wire			X41y84;
	wire			E51y84;
	wire			L51y84;
	wire			S51y84;
	wire			Z51y84;
	wire			G61y84;
	wire			N61y84;
	wire			U61y84;
	wire			B71y84;
	wire			I71y84;
	wire			P71y84;
	wire			W71y84;
	wire			D81y84;
	wire			K81y84;
	wire			R81y84;
	wire			Y81y84;
	wire			F91y84;
	wire			M91y84;
	wire			T91y84;
	wire			Aa1y84;
	wire			Ha1y84;
	wire			Oa1y84;
	wire			Va1y84;
	wire			Cb1y84;
	wire			Jb1y84;
	wire			Qb1y84;
	wire			Xb1y84;
	wire			Ec1y84;
	wire			Lc1y84;
	wire			Sc1y84;
	wire			Zc1y84;
	wire			Gd1y84;
	wire			Nd1y84;
	wire			Ud1y84;
	wire			Be1y84;
	wire			Ie1y84;
	wire			Pe1y84;
	wire			We1y84;
	wire			Df1y84;
	wire			Kf1y84;
	wire			Rf1y84;
	wire			Yf1y84;
	wire			Fg1y84;
	wire			Mg1y84;
	wire			Tg1y84;
	wire			Ah1y84;
	wire			Hh1y84;
	wire			Oh1y84;
	wire			Vh1y84;
	wire			Ci1y84;
	wire			Ji1y84;
	wire			Qi1y84;
	wire			Xi1y84;
	wire			Ej1y84;
	wire			Lj1y84;
	wire			Sj1y84;
	wire			Zj1y84;
	wire			Gk1y84;
	wire			Nk1y84;
	wire			Uk1y84;
	wire			Bl1y84;
	wire			Il1y84;
	wire			Pl1y84;
	wire			Wl1y84;
	wire			Dm1y84;
	wire			Km1y84;
	wire			Rm1y84;
	wire			Ym1y84;
	wire			Fn1y84;
	wire			Mn1y84;
	wire			Tn1y84;
	wire			Ao1y84;
	wire			Ho1y84;
	wire			Oo1y84;
	wire			Vo1y84;
	wire			Cp1y84;
	wire			Jp1y84;
	wire			Qp1y84;
	wire			Xp1y84;
	wire			Eq1y84;
	wire			Lq1y84;
	wire			Sq1y84;
	wire			Zq1y84;
	wire			Gr1y84;
	wire			Nr1y84;
	wire			Ur1y84;
	wire			Bs1y84;
	wire			Is1y84;
	wire			Ps1y84;
	wire			Ws1y84;
	wire			Dt1y84;
	wire			Kt1y84;
	wire			Rt1y84;
	wire			Yt1y84;
	wire			Fu1y84;
	wire			Mu1y84;
	wire			Tu1y84;
	wire			Av1y84;
	wire			Hv1y84;
	wire			Ov1y84;
	wire			Vv1y84;
	wire			Cw1y84;
	wire			Jw1y84;
	wire			Qw1y84;
	wire			Xw1y84;
	wire			Ex1y84;
	wire			Lx1y84;
	wire			Sx1y84;
	wire			Zx1y84;
	wire			Gy1y84;
	wire			Ny1y84;
	wire			Uy1y84;
	wire			Bz1y84;
	wire			Iz1y84;
	wire			Pz1y84;
	wire			Wz1y84;
	wire			D02y84;
	wire			K02y84;
	wire			R02y84;
	wire			Y02y84;
	wire			F12y84;
	wire			M12y84;
	wire			T12y84;
	wire			A22y84;
	wire			H22y84;
	wire			O22y84;
	wire			V22y84;
	wire			C32y84;
	wire			J32y84;
	wire			Q32y84;
	wire			X32y84;
	wire			E42y84;
	wire			L42y84;
	wire			S42y84;
	wire			Z42y84;
	wire			G52y84;
	wire			N52y84;
	wire			U52y84;
	wire			B62y84;
	wire			I62y84;
	wire			P62y84;
	wire			W62y84;
	wire			D72y84;
	wire			K72y84;
	wire			R72y84;
	wire			Y72y84;
	wire			F82y84;
	wire			M82y84;
	wire			T82y84;
	wire			A92y84;
	wire			H92y84;
	wire			O92y84;
	wire			V92y84;
	wire			Ca2y84;
	wire			Ja2y84;
	wire			Qa2y84;
	wire			Xa2y84;
	wire			Eb2y84;
	wire			Lb2y84;
	wire			Sb2y84;
	wire			Zb2y84;
	wire			Gc2y84;
	wire			Nc2y84;
	wire			Uc2y84;
	wire			Bd2y84;
	wire			Id2y84;
	wire			Pd2y84;
	wire			Wd2y84;
	wire			De2y84;
	wire			Mi42a4;
	wire			Ti42a4;
	wire			Aj42a4;
	wire			Hj42a4;
	wire			Oj42a4;
	wire			Vj42a4;
	wire			Ck42a4;
	wire			Jk42a4;
	wire			Qk42a4;
	wire			Xk42a4;
	wire			El42a4;
	wire			Ll42a4;
	wire			Sl42a4;
	wire			Zl42a4;
	wire			Gm42a4;
	wire			Nm42a4;
	wire			Um42a4;
	wire			Bn42a4;
	wire			In42a4;
	wire			Pn42a4;
	wire			Wn42a4;
	wire			Do42a4;
	wire			Ko42a4;
	wire			Ro42a4;
	wire			Yo42a4;
	wire			Fp42a4;
	wire			Mp42a4;
	wire			Tp42a4;
	wire			Aq42a4;
	wire			Hq42a4;
	wire			Oq42a4;
	wire			Vq42a4;
	wire			Cr42a4;
	wire			Jr42a4;
	wire			Qr42a4;
	wire			Xr42a4;
	wire			Es42a4;
	wire			Ls42a4;
	wire			Ss42a4;
	wire			Zs42a4;
	wire			Gt42a4;
	wire			Nt42a4;
	wire			Ut42a4;
	wire			Bu42a4;
	wire			Iu42a4;
	wire			Pu42a4;
	wire			Wu42a4;
	wire			Dv42a4;
	wire			Kv42a4;
	wire			Rv42a4;
	wire			Yv42a4;
	wire			Fw42a4;
	wire			Mw42a4;
	wire			Tw42a4;
	wire			Ax42a4;
	wire			Hx42a4;
	wire			Ox42a4;
	wire			Vx42a4;
	wire			Cy42a4;
	wire			Jy42a4;
	wire			Qy42a4;
	wire			Xy42a4;
	wire			Ez42a4;
	wire			Lz42a4;
	wire			Sz42a4;
	wire			Zz42a4;
	wire			G052a4;
	wire			N052a4;
	wire			U052a4;
	wire			B152a4;
	wire			I152a4;
	wire			P152a4;
	wire			W152a4;
	wire			D252a4;
	wire			K252a4;
	wire			R252a4;
	wire			Y252a4;
	wire			F352a4;
	wire			M352a4;
	wire			T352a4;
	wire			A452a4;
	wire			H452a4;
	wire			O452a4;
	wire			V452a4;
	wire			C552a4;
	wire			J552a4;
	wire			Q552a4;
	wire			X552a4;
	wire			E652a4;
	wire			L652a4;
	wire			S652a4;
	wire			Z652a4;
	wire			G752a4;
	wire			N752a4;
	wire			U752a4;
	wire			B852a4;
	wire			I852a4;
	wire			P852a4;
	wire			W852a4;
	wire			D952a4;
	wire			K952a4;
	wire			R952a4;
	wire			Y952a4;
	wire			Fa52a4;
	wire			Ma52a4;
	wire			Ta52a4;
	wire			Ab52a4;
	wire			Hb52a4;
	wire			Ob52a4;
	wire			Vb52a4;
	wire			Cc52a4;
	wire			Jc52a4;
	wire			Qc52a4;
	wire			Xc52a4;
	wire			Ed52a4;
	wire			Ld52a4;
	wire			Sd52a4;
	wire			Zd52a4;
	wire			Ge52a4;
	wire			Ne52a4;
	wire			Ue52a4;
	wire			Bf52a4;
	wire			If52a4;
	wire			Pf52a4;
	wire			Wf52a4;
	wire			Dg52a4;
	wire			Kg52a4;
	wire			Rg52a4;
	wire			Yg52a4;
	wire			Fh52a4;
	wire			Mh52a4;
	wire			Th52a4;
	wire			Ai52a4;
	wire			Hi52a4;
	wire			Oi52a4;
	wire			Vi52a4;
	wire			Cj52a4;
	wire			Jj52a4;
	wire			Qj52a4;
	wire			Xj52a4;
	wire			Ek52a4;
	wire			Lk52a4;
	wire			Sk52a4;
	wire			Zk52a4;
	wire			Gl52a4;
	wire			Nl52a4;
	wire			Ul52a4;
	wire			Bm52a4;
	wire			Im52a4;
	wire			Pm52a4;
	wire			Wm52a4;
	wire			Dn52a4;
	wire			Kn52a4;
	wire			Rn52a4;
	wire			Yn52a4;
	wire			Fo52a4;
	wire			Mo52a4;
	wire			To52a4;
	wire			Ap52a4;
	wire			Hp52a4;
	wire			Op52a4;
	wire			Vp52a4;
	wire			Cq52a4;
	wire			Jq52a4;
	wire			Qq52a4;
	wire			Xq52a4;
	wire			Er52a4;
	wire			Lr52a4;
	wire			Sr52a4;
	wire			Zr52a4;
	wire			Gs52a4;
	wire			Ns52a4;
	wire			Us52a4;
	wire			Bt52a4;
	wire			It52a4;
	wire			Pt52a4;
	wire			Wt52a4;
	wire			Du52a4;
	wire			Ku52a4;
	wire			Ru52a4;
	wire			Yu52a4;
	wire			Fv52a4;
	wire			Mv52a4;
	wire			Tv52a4;
	wire			Aw52a4;
	wire			Hw52a4;
	wire			Ow52a4;
	wire			Vw52a4;
	wire			Cx52a4;
	wire			Jx52a4;
	wire			Qx52a4;
	wire			Xx52a4;
	wire			Ey52a4;
	wire			Ly52a4;
	wire			Sy52a4;
	wire			Zy52a4;
	wire			Gz52a4;
	wire			Nz52a4;
	wire			Uz52a4;
	wire			B062a4;
	wire			I062a4;
	wire			P062a4;
	wire			W062a4;
	wire			D162a4;
	wire			K162a4;
	wire			R162a4;
	wire			Y162a4;
	wire			F262a4;
	wire			M262a4;
	wire			T262a4;
	wire			A362a4;
	wire			H362a4;
	wire			O362a4;
	wire			V362a4;
	wire			C462a4;
	wire			J462a4;
	wire			Q462a4;
	wire			X462a4;
	wire			E562a4;
	wire			L562a4;
	wire			S562a4;
	wire			Z562a4;
	wire			G662a4;
	wire			N662a4;
	wire			U662a4;
	wire			B762a4;
	wire			I762a4;
	wire			P762a4;
	wire			W762a4;
	wire			D862a4;
	wire			K862a4;
	wire			R862a4;
	wire			Y862a4;
	wire			F962a4;
	wire			M962a4;
	wire			T962a4;
	wire			Aa62a4;
	wire			Ha62a4;
	wire			Oa62a4;
	wire			Va62a4;
	wire			Cb62a4;
	wire			Jb62a4;
	wire			Qb62a4;
	wire			Xb62a4;
	wire			Ec62a4;
	wire			Lc62a4;
	wire			Sc62a4;
	wire			Zc62a4;
	wire			Gd62a4;
	wire			Nd62a4;
	wire			Ud62a4;
	wire			Be62a4;
	wire			Ie62a4;
	wire			Pe62a4;
	wire			We62a4;
	wire			Df62a4;
	wire			Kf62a4;
	wire			Rf62a4;
	wire			Yf62a4;
	wire			Fg62a4;
	wire			Mg62a4;
	wire			Tg62a4;
	wire			Ah62a4;
	wire			Hh62a4;
	wire			Oh62a4;
	wire			Vh62a4;
	wire			Ci62a4;
	wire			Ji62a4;
	wire			Qi62a4;
	wire			Xi62a4;
	wire			Ej62a4;
	wire			Lj62a4;
	wire			Sj62a4;
	wire			Zj62a4;
	wire			Gk62a4;
	wire			Nk62a4;
	wire			Uk62a4;
	wire			Bl62a4;
	wire			Il62a4;
	wire			Pl62a4;
	wire			Wl62a4;
	wire			Dm62a4;
	wire			Km62a4;
	wire			Rm62a4;
	wire			Ym62a4;
	wire			Fn62a4;
	wire			Mn62a4;
	wire			Tn62a4;
	wire			Ao62a4;
	wire			Ho62a4;
	wire			Oo62a4;
	wire			Vo62a4;
	wire			Cp62a4;
	wire			Jp62a4;
	wire			Qp62a4;
	wire			Xp62a4;
	wire			Eq62a4;
	wire			Lq62a4;
	wire			Sq62a4;
	wire			Zq62a4;
	wire			Gr62a4;
	wire			Nr62a4;
	wire			Ur62a4;
	wire			Bs62a4;
	wire			Is62a4;
	wire			Ps62a4;
	wire			Ws62a4;
	wire			Dt62a4;
	wire			Kt62a4;
	wire			Rt62a4;
	wire			Yt62a4;
	wire			Fu62a4;
	wire			Mu62a4;
	wire			Tu62a4;
	wire			Av62a4;
	wire			Hv62a4;
	wire			Ov62a4;
	wire			Vv62a4;
	wire			Cw62a4;
	wire			Jw62a4;
	wire			Qw62a4;
	wire			Xw62a4;
	wire			Ex62a4;
	wire			Lx62a4;
	wire			Sx62a4;
	wire			Zx62a4;
	wire			Gy62a4;
	wire			Ny62a4;
	wire			Uy62a4;
	wire			Bz62a4;
	wire			Iz62a4;
	wire			Pz62a4;
	wire			Wz62a4;
	wire			D072a4;
	wire			K072a4;
	wire			R072a4;
	wire			Y072a4;
	wire			F172a4;
	wire			M172a4;
	wire			T172a4;
	wire			A272a4;
	wire			H272a4;
	wire			O272a4;
	wire			V272a4;
	wire			C372a4;
	wire			J372a4;
	wire			Q372a4;
	wire			X372a4;
	wire			E472a4;
	wire			L472a4;
	wire			S472a4;
	wire			Z472a4;
	wire			G572a4;
	wire			N572a4;
	wire			U572a4;
	wire			B672a4;
	wire			I672a4;
	wire			P672a4;
	wire			W672a4;
	wire			D772a4;
	wire			K772a4;
	wire			R772a4;
	wire			Y772a4;
	wire			F872a4;
	wire			M872a4;
	wire			T872a4;
	wire			A972a4;
	wire			H972a4;
	wire			O972a4;
	wire			V972a4;
	wire			Ca72a4;
	wire			Ja72a4;
	wire			Qa72a4;
	wire			Xa72a4;
	wire			Eb72a4;
	wire			Lb72a4;
	wire			Sb72a4;
	wire			Zb72a4;
	wire			Gc72a4;
	wire			Nc72a4;
	wire			Uc72a4;
	wire			Bd72a4;
	wire			Id72a4;
	wire			Pd72a4;
	wire			Wd72a4;
	wire			De72a4;
	wire			Ke72a4;
	wire			Re72a4;
	wire			Ye72a4;
	wire			Ff72a4;
	wire			Mf72a4;
	wire			Tf72a4;
	wire			Ag72a4;
	wire			Hg72a4;
	wire			Og72a4;
	wire			Vg72a4;
	wire			Ch72a4;
	wire			Jh72a4;
	wire			Qh72a4;
	wire			Xh72a4;
	wire			Ei72a4;
	wire			Li72a4;
	wire			Si72a4;
	wire			Zi72a4;
	wire			Gj72a4;
	wire			Nj72a4;
	wire			Uj72a4;
	wire			Bk72a4;
	wire			Ik72a4;
	wire			Pk72a4;
	wire			Wk72a4;
	wire			Dl72a4;
	wire			Kl72a4;
	wire			Rl72a4;
	wire			Yl72a4;
	wire			Fm72a4;
	wire			Mm72a4;
	wire			Tm72a4;
	wire			An72a4;
	wire			Hn72a4;
	wire			On72a4;
	wire			Vn72a4;
	wire			Co72a4;
	wire			Jo72a4;
	wire			Qo72a4;
	wire			Xo72a4;
	wire			Ep72a4;
	wire			Lp72a4;
	wire			Sp72a4;
	wire			Zp72a4;
	wire			Gq72a4;
	wire			Nq72a4;
	wire			Uq72a4;
	wire			Br72a4;
	wire			Ir72a4;
	wire			Pr72a4;
	wire			Wr72a4;
	wire			Ds72a4;
	wire			Ks72a4;
	wire			Rs72a4;
	wire			Ys72a4;
	wire			Ft72a4;
	wire			Mt72a4;
	wire			Tt72a4;
	wire			Au72a4;
	wire			Hu72a4;
	wire			Ou72a4;
	wire			Vu72a4;
	wire			Cv72a4;
	wire			Jv72a4;
	wire			Qv72a4;
	wire			Xv72a4;
	wire			Ew72a4;
	wire			Lw72a4;
	wire			Sw72a4;
	wire			Zw72a4;
	wire			Gx72a4;
	wire			Nx72a4;
	wire			Ux72a4;
	wire			By72a4;
	wire			Iy72a4;
	wire			Py72a4;
	wire			Wy72a4;
	wire			Dz72a4;
	wire			Kz72a4;
	wire			Rz72a4;
	wire			Yz72a4;
	wire			F082a4;
	wire			M082a4;
	wire			T082a4;
	wire			A182a4;
	wire			H182a4;
	wire			O182a4;
	wire			V182a4;
	wire			C282a4;
	wire			J282a4;
	wire			Q282a4;
	wire			X282a4;
	wire			E382a4;
	wire			L382a4;
	wire			S382a4;
	wire			Z382a4;
	wire			G482a4;
	wire			N482a4;
	wire			U482a4;
	wire			B582a4;
	wire			I582a4;
	wire			P582a4;
	wire			W582a4;
	wire			D682a4;
	wire			K682a4;
	wire			R682a4;
	wire			Y682a4;
	wire			F782a4;
	wire			M782a4;
	wire			T782a4;
	wire			A882a4;
	wire			H882a4;
	wire			O882a4;
	wire			V882a4;
	wire			C982a4;
	wire			J982a4;
	wire			Q982a4;
	wire			X982a4;
	wire			Ea82a4;
	wire			La82a4;
	wire			Sa82a4;
	wire			Za82a4;
	wire			Gb82a4;
	wire			Nb82a4;
	wire			Ub82a4;
	wire			Bc82a4;
	wire			Ic82a4;
	wire			Pc82a4;
	wire			Wc82a4;
	wire			Dd82a4;
	wire			Kd82a4;
	wire			Rd82a4;
	wire			Yd82a4;
	wire			Fe82a4;
	wire			Me82a4;
	wire			Te82a4;
	wire			Af82a4;
	wire			Hf82a4;
	wire			Of82a4;
	wire			Vf82a4;
	wire			Cg82a4;
	wire			Jg82a4;
	wire			Qg82a4;
	wire			Xg82a4;
	wire			Eh82a4;
	wire			Lh82a4;
	wire			Sh82a4;
	wire			Zh82a4;
	wire			Gi82a4;
	wire			Ni82a4;
	wire			Ui82a4;
	wire			Bj82a4;
	wire			Ij82a4;
	wire			Pj82a4;
	wire			Wj82a4;
	wire			Dk82a4;
	wire			Kk82a4;
	wire			Rk82a4;
	wire			Yk82a4;
	wire			Fl82a4;
	wire			Ml82a4;
	wire			Tl82a4;
	wire			Am82a4;
	wire			Hm82a4;
	wire			Om82a4;
	wire			Vm82a4;
	wire			Cn82a4;
	wire			Jn82a4;
	wire			Qn82a4;
	wire			Xn82a4;
	wire			Eo82a4;
	wire			Lo82a4;
	wire			So82a4;
	wire			Zo82a4;
	wire			Gp82a4;
	wire			Np82a4;
	wire			Up82a4;
	wire			Bq82a4;
	wire			Iq82a4;
	wire			Pq82a4;
	wire			Wq82a4;
	wire			Dr82a4;
	wire			Kr82a4;
	wire			Rr82a4;
	wire			Yr82a4;
	wire			Fs82a4;
	wire			Ms82a4;
	wire			Ts82a4;
	wire			At82a4;
	wire			Ht82a4;
	wire			Ot82a4;
	wire			Vt82a4;
	wire			Cu82a4;
	wire			Ju82a4;
	wire			Qu82a4;
	wire			Xu82a4;
	wire			Ev82a4;
	wire			Lv82a4;
	wire			Sv82a4;
	wire			Zv82a4;
	wire			Gw82a4;
	wire			Nw82a4;
	wire			Uw82a4;
	wire			Bx82a4;
	wire			Ix82a4;
	wire			Px82a4;
	wire			Wx82a4;
	wire			Dy82a4;
	wire			Ky82a4;
	wire			Ry82a4;
	wire			Yy82a4;
	wire			Fz82a4;
	wire			Mz82a4;
	wire			Tz82a4;
	wire			A092a4;
	wire			H092a4;
	wire			O092a4;
	wire			V092a4;
	wire			C192a4;
	wire			J192a4;
	wire			Q192a4;
	wire			X192a4;
	wire			E292a4;
	wire			L292a4;
	wire			S292a4;
	wire			Z292a4;
	wire			G392a4;
	wire			N392a4;
	wire			U392a4;
	wire			B492a4;
	wire			I492a4;
	wire			P492a4;
	wire			W492a4;
	wire			D592a4;
	wire			K592a4;
	wire			R592a4;
	wire			Y592a4;
	wire			F692a4;
	wire			M692a4;
	wire			T692a4;
	wire			A792a4;
	wire			H792a4;
	wire			O792a4;
	wire			V792a4;
	wire			C892a4;
	wire			J892a4;
	wire			Q892a4;
	wire			X892a4;
	wire			E992a4;
	wire			L992a4;
	wire			S992a4;
	wire			Z992a4;
	wire			Ga92a4;
	wire			Na92a4;
	wire			Ua92a4;
	wire			Bb92a4;
	wire			Ib92a4;
	wire			Pb92a4;
	wire			Wb92a4;
	wire			Dc92a4;
	wire			Kc92a4;
	wire			Rc92a4;
	wire			Yc92a4;
	wire			Fd92a4;
	wire			Md92a4;
	wire			Td92a4;
	wire			Ae92a4;
	wire			He92a4;
	wire			Oe92a4;
	wire			Ve92a4;
	wire			Cf92a4;
	wire			Jf92a4;
	wire			Qf92a4;
	wire			Xf92a4;
	wire			Eg92a4;
	wire			Lg92a4;
	wire			Sg92a4;
	wire			Zg92a4;
	wire			Gh92a4;
	wire			Nh92a4;
	wire			Uh92a4;
	wire			Bi92a4;
	wire			Ii92a4;
	wire			Pi92a4;
	wire			Wi92a4;
	wire			Dj92a4;
	wire			Kj92a4;
	wire			Rj92a4;
	wire			Yj92a4;
	wire			Fk92a4;
	wire			Mk92a4;
	wire			Tk92a4;
	wire			Al92a4;
	wire			Hl92a4;
	wire			Ol92a4;
	wire			Vl92a4;
	wire			Cm92a4;
	wire			Jm92a4;
	wire			Qm92a4;
	wire			Xm92a4;
	wire			En92a4;
	wire			Ln92a4;
	wire			Sn92a4;
	wire			Zn92a4;
	wire			Go92a4;
	wire			No92a4;
	wire			Uo92a4;
	wire			Bp92a4;
	wire			Ip92a4;
	wire			Pp92a4;
	wire			Wp92a4;
	wire			Dq92a4;
	wire			Kq92a4;
	wire			Rq92a4;
	wire			Yq92a4;
	wire			Fr92a4;
	wire			Mr92a4;
	wire			Tr92a4;
	wire			As92a4;
	wire			Hs92a4;
	wire			Os92a4;
	wire			Vs92a4;
	wire			Ct92a4;
	wire			Jt92a4;
	wire			Qt92a4;
	wire			Xt92a4;
	wire			Eu92a4;
	wire			Lu92a4;
	wire			Su92a4;
	wire			Zu92a4;
	wire			Gv92a4;
	wire			Nv92a4;
	wire			Uv92a4;
	wire			Bw92a4;
	wire			Iw92a4;
	wire			Pw92a4;
	wire			Ww92a4;
	wire			Dx92a4;
	wire			Kx92a4;
	wire			Rx92a4;
	wire			Yx92a4;
	wire			Fy92a4;
	wire			My92a4;
	wire			Ty92a4;
	wire			Az92a4;
	wire			Hz92a4;
	wire			Oz92a4;
	wire			Vz92a4;
	wire			C0a2a4;
	wire			J0a2a4;
	wire			Q0a2a4;
	wire			X0a2a4;
	wire			E1a2a4;
	wire			L1a2a4;
	wire			S1a2a4;
	wire			Z1a2a4;
	wire			G2a2a4;
	wire			N2a2a4;
	wire			U2a2a4;
	wire			B3a2a4;
	wire			I3a2a4;
	wire			P3a2a4;
	wire			W3a2a4;
	wire			D4a2a4;
	wire			K4a2a4;
	wire			R4a2a4;
	wire			Y4a2a4;
	wire			F5a2a4;
	wire			M5a2a4;
	wire			T5a2a4;
	wire			A6a2a4;
	wire			H6a2a4;
	wire			O6a2a4;
	wire			V6a2a4;
	wire			C7a2a4;
	wire			J7a2a4;
	wire			Q7a2a4;
	wire			X7a2a4;
	wire			E8a2a4;
	wire			L8a2a4;
	wire			S8a2a4;
	wire			Z8a2a4;
	wire			G9a2a4;
	wire			N9a2a4;
	wire			U9a2a4;
	wire			Baa2a4;
	wire			Iaa2a4;
	wire			Paa2a4;
	wire			Waa2a4;
	wire			Dba2a4;
	wire			Kba2a4;
	wire			Rba2a4;
	wire			Yba2a4;
	wire			Fca2a4;
	wire			Mca2a4;
	wire			Tca2a4;
	wire			Ada2a4;
	wire			Hda2a4;
	wire			Oda2a4;
	wire			Vda2a4;
	wire			Cea2a4;
	wire			Jea2a4;
	wire			Qea2a4;
	wire			Xea2a4;
	wire			Efa2a4;
	wire			Lfa2a4;
	wire			Sfa2a4;
	wire			Zfa2a4;
	wire			Gga2a4;
	wire			Nga2a4;
	wire			Uga2a4;
	wire			Bha2a4;
	wire			Iha2a4;
	wire			Pha2a4;
	wire			Wha2a4;
	wire			Dia2a4;
	wire			Kia2a4;
	wire			Ria2a4;
	wire			Yia2a4;
	wire			Fja2a4;
	wire			Mja2a4;
	wire			Tja2a4;
	wire			Aka2a4;
	wire			Hka2a4;
	wire			Oka2a4;
	wire			Vka2a4;
	wire			Cla2a4;
	wire			Jla2a4;
	wire			Qla2a4;
	wire			Xla2a4;
	wire			Ema2a4;
	wire			Lma2a4;
	wire			Sma2a4;
	wire			Zma2a4;
	wire			Gna2a4;
	wire			Nna2a4;
	wire			Una2a4;
	wire			Boa2a4;
	wire			Ioa2a4;
	wire			Poa2a4;
	wire			Woa2a4;
	wire			Dpa2a4;
	wire			Kpa2a4;
	wire			Rpa2a4;
	wire			Ypa2a4;
	wire			Fqa2a4;
	wire			Mqa2a4;
	wire			Tqa2a4;
	wire			Ara2a4;
	wire			Hra2a4;
	wire			Ora2a4;
	wire			Vra2a4;
	wire			Csa2a4;
	wire			Jsa2a4;
	wire			Qsa2a4;
	wire			Xsa2a4;
	wire			Eta2a4;
	wire			Lta2a4;
	wire			Sta2a4;
	wire			Zta2a4;
	wire			Gua2a4;
	wire			Nua2a4;
	wire			Uua2a4;
	wire			Bva2a4;
	wire			Iva2a4;
	wire			Pva2a4;
	wire			Wva2a4;
	wire			Dwa2a4;
	wire			Kwa2a4;
	wire			Rwa2a4;
	wire			Ywa2a4;
	wire			Fxa2a4;
	wire			Mxa2a4;
	wire			Txa2a4;
	wire			Aya2a4;
	wire			Hya2a4;
	wire			Oya2a4;
	wire			Vya2a4;
	wire			Cza2a4;
	wire			Jza2a4;
	wire			Qza2a4;
	wire			Xza2a4;
	wire			E0b2a4;
	wire			L0b2a4;
	wire			S0b2a4;
	wire			Z0b2a4;
	wire			G1b2a4;
	wire			N1b2a4;
	wire			U1b2a4;
	wire			B2b2a4;
	wire			I2b2a4;
	wire			P2b2a4;
	wire			W2b2a4;
	wire			D3b2a4;
	wire			K3b2a4;
	wire			R3b2a4;
	wire			Y3b2a4;
	wire			F4b2a4;
	wire			M4b2a4;
	wire			T4b2a4;
	wire			A5b2a4;
	wire			H5b2a4;
	wire			O5b2a4;
	wire			V5b2a4;
	wire			C6b2a4;
	wire			J6b2a4;
	wire			Q6b2a4;
	wire			X6b2a4;
	wire			E7b2a4;
	wire			L7b2a4;
	wire			S7b2a4;
	wire			Z7b2a4;
	wire			G8b2a4;
	wire			N8b2a4;
	wire			U8b2a4;
	wire			B9b2a4;
	wire			I9b2a4;
	wire			P9b2a4;
	wire			W9b2a4;
	wire			Dab2a4;
	wire			Kab2a4;
	wire			Rab2a4;
	wire			Yab2a4;
	wire			Fbb2a4;
	wire			Mbb2a4;
	wire			Tbb2a4;
	wire			Acb2a4;
	wire			Hcb2a4;
	wire			Ocb2a4;
	wire			Vcb2a4;
	wire			Cdb2a4;
	wire			Jdb2a4;
	wire			Qdb2a4;
	wire			Xdb2a4;
	wire			Eeb2a4;
	wire			Leb2a4;
	wire			Seb2a4;
	wire			Zeb2a4;
	wire			Gfb2a4;
	wire			Nfb2a4;
	wire			Ufb2a4;
	wire			Bgb2a4;
	wire			Igb2a4;
	wire			Pgb2a4;
	wire			Wgb2a4;
	wire			Dhb2a4;
	wire			Khb2a4;
	wire			Rhb2a4;
	wire			Yhb2a4;
	wire			Fib2a4;
	wire			Mib2a4;
	wire			Tib2a4;
	wire			Ajb2a4;
	wire			Hjb2a4;
	wire			Ojb2a4;
	wire			Vjb2a4;
	wire			Ckb2a4;
	wire			Jkb2a4;
	wire			Qkb2a4;
	wire			Xkb2a4;
	wire			Elb2a4;
	wire			Llb2a4;
	wire			Slb2a4;
	wire			Zlb2a4;
	wire			Gmb2a4;
	wire			Nmb2a4;
	wire			Umb2a4;
	wire			Bnb2a4;
	wire			Inb2a4;
	wire			Pnb2a4;
	wire			Wnb2a4;
	wire			Dob2a4;
	wire			Kob2a4;
	wire			Rob2a4;
	wire			Yob2a4;
	wire			Fpb2a4;
	wire			Mpb2a4;
	wire			Tpb2a4;
	wire			Aqb2a4;
	wire			Hqb2a4;
	wire			Oqb2a4;
	wire			Vqb2a4;
	wire			Crb2a4;
	wire			Jrb2a4;
	wire			Qrb2a4;
	wire			Xrb2a4;
	wire			Esb2a4;
	wire			Lsb2a4;
	wire			Ssb2a4;
	wire			Zsb2a4;
	wire			Gtb2a4;
	wire			Ntb2a4;
	wire			Utb2a4;
	wire			Bub2a4;
	wire			Iub2a4;
	wire			Pub2a4;
	wire			Wub2a4;
	wire			Dvb2a4;
	wire			Kvb2a4;
	wire			Rvb2a4;
	wire			Yvb2a4;
	wire			Fwb2a4;
	wire			Mwb2a4;
	wire			Twb2a4;
	wire			Axb2a4;
	wire			Hxb2a4;
	wire			Oxb2a4;
	wire			Vxb2a4;
	wire			Cyb2a4;
	wire			Jyb2a4;
	wire			Qyb2a4;
	wire			Xyb2a4;
	wire			Ezb2a4;
	wire			Lzb2a4;
	wire			Szb2a4;
	wire			Zzb2a4;
	wire			G0c2a4;
	wire			N0c2a4;
	wire			U0c2a4;
	wire			B1c2a4;
	wire			I1c2a4;
	wire			P1c2a4;
	wire			W1c2a4;
	wire			D2c2a4;
	wire			K2c2a4;
	wire			R2c2a4;
	wire			Y2c2a4;
	wire			F3c2a4;
	wire			M3c2a4;
	wire			T3c2a4;
	wire			A4c2a4;
	wire			H4c2a4;
	wire			O4c2a4;
	wire			V4c2a4;
	wire			C5c2a4;
	wire			J5c2a4;
	wire			Q5c2a4;
	wire			X5c2a4;
	wire			E6c2a4;
	wire			L6c2a4;
	wire			S6c2a4;
	wire			Z6c2a4;
	wire			G7c2a4;
	wire			N7c2a4;
	wire			U7c2a4;
	wire			B8c2a4;
	wire			I8c2a4;
	wire			P8c2a4;
	wire			W8c2a4;
	wire			D9c2a4;
	wire			K9c2a4;
	wire			R9c2a4;
	wire			Y9c2a4;
	wire			Fac2a4;
	wire			Mac2a4;
	wire			Tac2a4;
	wire			Abc2a4;
	wire			Hbc2a4;
	wire			Obc2a4;
	wire			Vbc2a4;
	wire			Ccc2a4;
	wire			Jcc2a4;
	wire			Qcc2a4;
	wire			Xcc2a4;
	wire			Edc2a4;
	wire			Ldc2a4;
	wire			Sdc2a4;
	wire			Zdc2a4;
	wire			Gec2a4;
	wire			Nec2a4;
	wire			Uec2a4;
	wire			Bfc2a4;
	wire			Ifc2a4;
	wire			Pfc2a4;
	wire			Wfc2a4;
	wire			Dgc2a4;
	wire			Kgc2a4;
	wire			Rgc2a4;
	wire			Ygc2a4;
	wire			Fhc2a4;
	wire			Mhc2a4;
	wire			Thc2a4;
	wire			Aic2a4;
	wire			Hic2a4;
	wire			Oic2a4;
	wire			Vic2a4;
	wire			Cjc2a4;
	wire			Jjc2a4;
	wire			Qjc2a4;
	wire			Xjc2a4;
	wire			Ekc2a4;
	wire			Lkc2a4;
	wire			Skc2a4;
	wire			Zkc2a4;
	wire			Glc2a4;
	wire			Nlc2a4;
	wire			Ulc2a4;
	wire			Bmc2a4;
	wire			Imc2a4;
	wire			Pmc2a4;
	wire			Wmc2a4;
	wire			Dnc2a4;
	wire			Knc2a4;
	wire			Rnc2a4;
	wire			Ync2a4;
	wire			Foc2a4;
	wire			Moc2a4;
	wire			Toc2a4;
	wire			Apc2a4;
	wire			Hpc2a4;
	wire			Opc2a4;
	wire			Vpc2a4;
	wire			Cqc2a4;
	wire			Jqc2a4;
	wire			Qqc2a4;
	wire			Xqc2a4;
	wire			Erc2a4;
	wire			Lrc2a4;
	wire			Src2a4;
	wire			Zrc2a4;
	wire			Gsc2a4;
	wire			Nsc2a4;
	wire			Usc2a4;
	wire			Btc2a4;
	wire			Itc2a4;
	wire			Ptc2a4;
	wire			Wtc2a4;
	wire			Duc2a4;
	wire			Kuc2a4;
	wire			Ruc2a4;
	wire			Yuc2a4;
	wire			Fvc2a4;
	wire			Mvc2a4;
	wire			Tvc2a4;
	wire			Awc2a4;
	wire			Hwc2a4;
	wire			Owc2a4;
	wire			Vwc2a4;
	wire			Cxc2a4;
	wire			Jxc2a4;
	wire			Qxc2a4;
	wire			Xxc2a4;
	wire			Eyc2a4;
	wire			Lyc2a4;
	wire			Syc2a4;
	wire			Zyc2a4;
	wire			Gzc2a4;
	wire			Nzc2a4;
	wire			Uzc2a4;
	wire			B0d2a4;
	wire			I0d2a4;
	wire			P0d2a4;
	wire			W0d2a4;
	wire			D1d2a4;
	wire			K1d2a4;
	wire			R1d2a4;
	wire			Y1d2a4;
	wire			F2d2a4;
	wire			M2d2a4;
	wire			T2d2a4;
	wire			A3d2a4;
	wire			H3d2a4;
	wire			O3d2a4;
	wire			V3d2a4;
	wire			C4d2a4;
	wire			J4d2a4;
	wire			Q4d2a4;
	wire			X4d2a4;
	wire			E5d2a4;
	wire			L5d2a4;
	wire			S5d2a4;
	wire			Z5d2a4;
	wire			G6d2a4;
	wire			N6d2a4;
	wire			U6d2a4;
	wire			B7d2a4;
	wire			I7d2a4;
	wire			P7d2a4;
	wire			W7d2a4;
	wire			D8d2a4;
	wire			K8d2a4;
	wire			R8d2a4;
	wire			Y8d2a4;
	wire			F9d2a4;
	wire			M9d2a4;
	wire			T9d2a4;
	wire			Aad2a4;
	wire			Had2a4;
	wire			Oad2a4;
	wire			Vad2a4;
	wire			Cbd2a4;
	wire			Jbd2a4;
	wire			Qbd2a4;
	wire			Xbd2a4;
	wire			Ecd2a4;
	wire			Lcd2a4;
	wire			Scd2a4;
	wire			Zcd2a4;
	wire			Gdd2a4;
	wire			Ndd2a4;
	wire			Udd2a4;
	wire			Bed2a4;
	wire			Ied2a4;
	wire			Ped2a4;
	wire			Wed2a4;
	wire			Dfd2a4;
	wire			Kfd2a4;
	wire			Rfd2a4;
	wire			Yfd2a4;
	wire			Fgd2a4;
	wire			Mgd2a4;
	wire			Tgd2a4;
	wire			Ahd2a4;
	wire			Hhd2a4;
	wire			Ohd2a4;
	wire			Vhd2a4;
	wire			Cid2a4;
	wire			Jid2a4;
	wire			Qid2a4;
	wire			Xid2a4;
	wire			Ejd2a4;
	wire			Ljd2a4;
	wire			Sjd2a4;
	wire			Zjd2a4;
	wire			Gkd2a4;
	wire			Nkd2a4;
	wire			Ukd2a4;
	wire			Bld2a4;
	wire			Ild2a4;
	wire			Pld2a4;
	wire			Wld2a4;
	wire			Dmd2a4;
	wire			Kmd2a4;
	wire			Rmd2a4;
	wire			Ymd2a4;
	wire			Fnd2a4;
	wire			Mnd2a4;
	wire			Tnd2a4;
	wire			Aod2a4;
	wire			Hod2a4;
	wire			Ood2a4;
	wire			Vod2a4;
	wire			Cpd2a4;
	wire			Jpd2a4;
	wire			Qpd2a4;
	wire			Xpd2a4;
	wire			Eqd2a4;
	wire			Lqd2a4;
	wire			Sqd2a4;
	wire			Zqd2a4;
	wire			Grd2a4;
	wire			Nrd2a4;
	wire			Urd2a4;
	wire			Bsd2a4;
	wire			Isd2a4;
	wire			Psd2a4;
	wire			Wsd2a4;
	wire			Dtd2a4;
	wire			Ktd2a4;
	wire			Rtd2a4;
	wire			Ytd2a4;
	wire			Fud2a4;
	wire			Mud2a4;
	wire			Tud2a4;
	wire			Avd2a4;
	wire			Hvd2a4;
	wire			Ovd2a4;
	wire			Vvd2a4;
	wire			Cwd2a4;
	wire			Jwd2a4;
	wire			Qwd2a4;
	wire			Xwd2a4;
	wire			Exd2a4;
	wire			Lxd2a4;
	wire			Sxd2a4;
	wire			Zxd2a4;
	wire			Gyd2a4;
	wire			Nyd2a4;
	wire			Uyd2a4;
	wire			Bzd2a4;
	wire			Izd2a4;
	wire			Pzd2a4;
	wire			Wzd2a4;
	wire			D0e2a4;
	wire			K0e2a4;
	wire			R0e2a4;
	wire			Y0e2a4;
	wire			F1e2a4;
	wire			M1e2a4;
	wire			T1e2a4;
	wire			A2e2a4;
	wire			H2e2a4;
	wire			O2e2a4;
	wire			V2e2a4;
	wire			C3e2a4;
	wire			J3e2a4;
	wire			Q3e2a4;
	wire			X3e2a4;
	wire			E4e2a4;
	wire			L4e2a4;
	wire			S4e2a4;
	wire			Z4e2a4;
	wire			G5e2a4;
	wire			N5e2a4;
	wire			U5e2a4;
	wire			B6e2a4;
	wire			I6e2a4;
	wire			P6e2a4;
	wire			W6e2a4;
	wire			D7e2a4;
	wire			K7e2a4;
	wire			R7e2a4;
	wire			Y7e2a4;
	wire			F8e2a4;
	wire			M8e2a4;
	wire			T8e2a4;
	wire			A9e2a4;
	wire			H9e2a4;
	wire			O9e2a4;
	wire			V9e2a4;
	wire			Cae2a4;
	wire			Jae2a4;
	wire			Qae2a4;
	wire			Xae2a4;
	wire			Ebe2a4;
	wire			Lbe2a4;
	wire			Sbe2a4;
	wire			Zbe2a4;
	wire			Gce2a4;
	wire			Nce2a4;
	wire			Uce2a4;
	wire			Bde2a4;
	wire			Ide2a4;
	wire			Pde2a4;
	wire			Wde2a4;
	wire			Dee2a4;
	wire			Kee2a4;
	wire			Ree2a4;
	wire			Yee2a4;
	wire			Ffe2a4;
	wire			Mfe2a4;
	wire			Tfe2a4;
	wire			Age2a4;
	wire			Hge2a4;
	wire			Oge2a4;
	wire			Vge2a4;
	wire			Che2a4;
	wire			Jhe2a4;
	wire			Qhe2a4;
	wire			Xhe2a4;
	wire			Eie2a4;
	wire			Lie2a4;
	wire			Sie2a4;
	wire			Zie2a4;
	wire			Gje2a4;
	wire			Nje2a4;
	wire			Uje2a4;
	wire			Bke2a4;
	wire			Ike2a4;
	wire			Pke2a4;
	wire			Wke2a4;
	wire			Dle2a4;
	wire			Kle2a4;
	wire			Rle2a4;
	wire			Yle2a4;
	wire			Fme2a4;
	wire			Mme2a4;
	wire			Tme2a4;
	wire			Ane2a4;
	wire			Hne2a4;
	wire			One2a4;
	wire			Vne2a4;
	wire			Coe2a4;
	wire			Joe2a4;
	wire			Qoe2a4;
	wire			Xoe2a4;
	wire			Epe2a4;
	wire			Lpe2a4;
	wire			Spe2a4;
	wire			Zpe2a4;
	wire			Gqe2a4;
	wire			Nqe2a4;
	wire			Uqe2a4;
	wire			Bre2a4;
	wire			Ire2a4;
	wire			Pre2a4;
	wire			Wre2a4;
	wire			Dse2a4;
	wire			Kse2a4;
	wire			Rse2a4;
	wire			Yse2a4;
	wire			Fte2a4;
	wire			Mte2a4;
	wire			Tte2a4;
	wire			Aue2a4;
	wire			Hue2a4;
	wire			Oue2a4;
	wire			Vue2a4;
	wire			Cve2a4;
	wire			Jve2a4;
	wire			Qve2a4;
	wire			Xve2a4;
	wire			Ewe2a4;
	wire			Lwe2a4;
	wire			Swe2a4;
	wire			Zwe2a4;
	wire			Gxe2a4;
	wire			Nxe2a4;
	wire			Uxe2a4;
	wire			Bye2a4;
	wire			Iye2a4;
	wire			Pye2a4;
	wire			Wye2a4;
	wire			Dze2a4;
	wire			Kze2a4;
	wire			Rze2a4;
	wire			Yze2a4;
	wire			F0f2a4;
	wire			M0f2a4;
	wire			T0f2a4;
	wire			A1f2a4;
	wire			H1f2a4;
	wire			O1f2a4;
	wire			V1f2a4;
	wire			C2f2a4;
	wire			J2f2a4;
	wire			Q2f2a4;
	wire			X2f2a4;
	wire			E3f2a4;
	wire			L3f2a4;
	wire			S3f2a4;
	wire			Z3f2a4;
	wire			G4f2a4;
	wire			N4f2a4;
	wire			U4f2a4;
	wire			B5f2a4;
	wire			I5f2a4;
	wire			P5f2a4;
	wire			W5f2a4;
	wire			D6f2a4;
	wire			K6f2a4;
	wire			R6f2a4;
	wire			Y6f2a4;
	wire			F7f2a4;
	wire			M7f2a4;
	wire			T7f2a4;
	wire			A8f2a4;
	wire			H8f2a4;
	wire			O8f2a4;
	wire			V8f2a4;
	wire			C9f2a4;
	wire			J9f2a4;
	wire			Q9f2a4;
	wire			X9f2a4;
	wire			Eaf2a4;
	wire			Laf2a4;
	wire			Saf2a4;
	wire			Zaf2a4;
	wire			Gbf2a4;
	wire			Nbf2a4;
	wire			Ubf2a4;
	wire			Bcf2a4;
	wire			Icf2a4;
	wire			Pcf2a4;
	wire			Wcf2a4;
	wire			Ddf2a4;
	wire			Kdf2a4;
	wire			Rdf2a4;
	wire			Ydf2a4;
	wire			Fef2a4;
	wire			Mef2a4;
	wire			Tef2a4;
	wire			Aff2a4;
	wire			Hff2a4;
	wire			Off2a4;
	wire			Vff2a4;
	wire			Cgf2a4;
	wire			Jgf2a4;
	wire			Qgf2a4;
	wire			Xgf2a4;
	wire			Ehf2a4;
	wire			Lhf2a4;
	wire			Shf2a4;
	wire			Zhf2a4;
	wire			Gif2a4;
	wire			Nif2a4;
	wire			Uif2a4;
	wire			Bjf2a4;
	wire			Ijf2a4;
	wire			Pjf2a4;
	wire			Wjf2a4;
	wire			Dkf2a4;
	wire			Kkf2a4;
	wire			Rkf2a4;
	wire			Ykf2a4;
	wire			Flf2a4;
	wire			Mlf2a4;
	wire			Tlf2a4;
	wire			Amf2a4;
	wire			Hmf2a4;
	wire			Omf2a4;
	wire			Vmf2a4;
	wire			Cnf2a4;
	wire			Jnf2a4;
	wire			Qnf2a4;
	wire			Xnf2a4;
	wire			Eof2a4;
	wire			Lof2a4;
	wire			Sof2a4;
	wire			Zof2a4;
	wire			Gpf2a4;
	wire			Npf2a4;
	wire			Upf2a4;
	wire			Bqf2a4;
	wire			Iqf2a4;
	wire			Pqf2a4;
	wire			Wqf2a4;
	wire			Drf2a4;
	wire			Krf2a4;
	wire			Rrf2a4;
	wire			Yrf2a4;
	wire			Fsf2a4;
	wire			Msf2a4;
	wire			Tsf2a4;
	wire			Atf2a4;
	wire			Htf2a4;
	wire			Otf2a4;
	wire			Vtf2a4;
	wire			Cuf2a4;
	wire			Juf2a4;
	wire			Quf2a4;
	wire			Xuf2a4;
	wire			Evf2a4;
	wire			Lvf2a4;
	wire			Svf2a4;
	wire			Zvf2a4;
	wire			Gwf2a4;
	wire			Nwf2a4;
	wire			Uwf2a4;
	wire			Bxf2a4;
	wire			Ixf2a4;
	wire			Pxf2a4;
	wire			Wxf2a4;
	wire			Dyf2a4;
	wire			Kyf2a4;
	wire			Ryf2a4;
	wire			Yyf2a4;
	wire			Fzf2a4;
	wire			Mzf2a4;
	wire			Tzf2a4;
	wire			A0g2a4;
	wire			H0g2a4;
	wire			O0g2a4;
	wire			V0g2a4;
	wire			C1g2a4;
	wire			J1g2a4;
	wire			Q1g2a4;
	wire			X1g2a4;
	wire			E2g2a4;
	wire			L2g2a4;
	wire			S2g2a4;
	wire			Z2g2a4;
	wire			G3g2a4;
	wire			N3g2a4;
	wire			U3g2a4;
	wire			B4g2a4;
	wire			I4g2a4;
	wire			P4g2a4;
	wire			W4g2a4;
	wire			D5g2a4;
	wire			K5g2a4;
	wire			R5g2a4;
	wire			Y5g2a4;
	wire			F6g2a4;
	wire			M6g2a4;
	wire			T6g2a4;
	wire			A7g2a4;
	wire			H7g2a4;
	wire			O7g2a4;
	wire			V7g2a4;
	wire			C8g2a4;
	wire			J8g2a4;
	wire			Q8g2a4;
	wire			X8g2a4;
	wire			E9g2a4;
	wire			L9g2a4;
	wire			S9g2a4;
	wire			Z9g2a4;
	wire			Gag2a4;
	wire			Nag2a4;
	wire			Uag2a4;
	wire			Bbg2a4;
	wire			Ibg2a4;
	wire			Pbg2a4;
	wire			Wbg2a4;
	wire			Dcg2a4;
	wire			Kcg2a4;
	wire			Rcg2a4;
	wire			Ycg2a4;
	wire			Fdg2a4;
	wire			Mdg2a4;
	wire			Tdg2a4;
	wire			Aeg2a4;
	wire			Heg2a4;
	wire			Oeg2a4;
	wire			Veg2a4;
	wire			Cfg2a4;
	wire			Jfg2a4;
	wire			Qfg2a4;
	wire			Xfg2a4;
	wire			Egg2a4;
	wire			Lgg2a4;
	wire			Sgg2a4;
	wire			Zgg2a4;
	wire			Ghg2a4;
	wire			Nhg2a4;
	wire			Uhg2a4;
	wire			Big2a4;
	wire			Iig2a4;
	wire			Pig2a4;
	wire			Wig2a4;
	wire			Djg2a4;
	wire			Kjg2a4;
	wire			Rjg2a4;
	wire			Yjg2a4;
	wire			Fkg2a4;
	wire			Mkg2a4;
	wire			Tkg2a4;
	wire			Alg2a4;
	wire			Hlg2a4;
	wire			Olg2a4;
	wire			Vlg2a4;
	wire			Cmg2a4;
	wire			Jmg2a4;
	wire			Qmg2a4;
	wire			Xmg2a4;
	wire			Eng2a4;
	wire			Lng2a4;
	wire			Sng2a4;
	wire			Zng2a4;
	wire			Gog2a4;
	wire			Nog2a4;
	wire			Uog2a4;
	wire			Bpg2a4;
	wire			Ipg2a4;
	wire			Ppg2a4;
	wire			Wpg2a4;
	wire			Dqg2a4;
	wire			Kqg2a4;
	wire			Rqg2a4;
	wire			Yqg2a4;
	wire			Frg2a4;
	wire			Mrg2a4;
	wire			Trg2a4;
	wire			Asg2a4;
	wire			Hsg2a4;
	wire			Osg2a4;
	wire			Vsg2a4;
	wire			Ctg2a4;
	wire			Jtg2a4;
	wire			Qtg2a4;
	wire			Xtg2a4;
	wire			Eug2a4;
	wire			Lug2a4;
	wire			Sug2a4;
	wire			Zug2a4;
	wire			Gvg2a4;
	wire			Nvg2a4;
	wire			Uvg2a4;
	wire			Bwg2a4;
	wire			Iwg2a4;
	wire			Pwg2a4;
	wire			Wwg2a4;
	wire			Dxg2a4;
	wire			Kxg2a4;
	wire			Rxg2a4;
	wire			Yxg2a4;
	wire			Fyg2a4;
	wire			Myg2a4;
	wire			Tyg2a4;
	wire			Azg2a4;
	wire			Hzg2a4;
	wire			Ozg2a4;
	wire			Vzg2a4;
	wire			C0h2a4;
	wire			J0h2a4;
	wire			Q0h2a4;
	wire			X0h2a4;
	wire			E1h2a4;
	wire			L1h2a4;
	wire			S1h2a4;
	wire			Z1h2a4;
	wire			G2h2a4;
	wire			N2h2a4;
	wire			U2h2a4;
	wire			B3h2a4;
	wire			I3h2a4;
	wire			P3h2a4;
	wire			W3h2a4;
	wire			D4h2a4;
	wire			K4h2a4;
	wire			R4h2a4;
	wire			Y4h2a4;
	wire			F5h2a4;
	wire			M5h2a4;
	wire			T5h2a4;
	wire			A6h2a4;
	wire			H6h2a4;
	wire			O6h2a4;
	wire			V6h2a4;
	wire			C7h2a4;
	wire			J7h2a4;
	wire			Q7h2a4;
	wire			X7h2a4;
	wire			E8h2a4;
	wire			L8h2a4;
	wire			S8h2a4;
	wire			Z8h2a4;
	wire			G9h2a4;
	wire			N9h2a4;
	wire			U9h2a4;
	wire			Bah2a4;
	wire			Iah2a4;
	wire			Pah2a4;
	wire			Wah2a4;
	wire			Dbh2a4;
	wire			Kbh2a4;
	wire			Rbh2a4;
	wire			Ybh2a4;
	wire			Fch2a4;
	wire			Mch2a4;
	wire			Tch2a4;
	wire			Adh2a4;
	wire			Hdh2a4;
	wire			Odh2a4;
	wire			Vdh2a4;
	wire			Ceh2a4;
	wire			Jeh2a4;
	wire			Qeh2a4;
	wire			Xeh2a4;
	wire			Efh2a4;
	wire			Lfh2a4;
	wire			Sfh2a4;
	wire			Zfh2a4;
	wire			Ggh2a4;
	wire			Ngh2a4;
	wire			Ugh2a4;
	wire			Bhh2a4;
	wire			Ihh2a4;
	wire			Phh2a4;
	wire			Whh2a4;
	wire			Dih2a4;
	wire			Kih2a4;
	wire			Rih2a4;
	wire			Yih2a4;
	wire			Fjh2a4;
	wire			Mjh2a4;
	wire			Tjh2a4;
	wire			Akh2a4;
	wire			Hkh2a4;
	wire			Okh2a4;
	wire			Vkh2a4;
	wire			Clh2a4;
	wire			Jlh2a4;
	wire			Qlh2a4;
	wire			Xlh2a4;
	wire			Emh2a4;
	wire			Lmh2a4;
	wire			Smh2a4;
	wire			Zmh2a4;
	wire			Gnh2a4;
	wire			Nnh2a4;
	wire			Unh2a4;
	wire			Boh2a4;
	wire			Ioh2a4;
	wire			Poh2a4;
	wire			Woh2a4;
	wire			Dph2a4;
	wire			Kph2a4;
	wire			Rph2a4;
	wire			Yph2a4;
	wire			Fqh2a4;
	wire			Mqh2a4;
	wire			Tqh2a4;
	wire			Arh2a4;
	wire			Hrh2a4;
	wire			Orh2a4;
	wire			Vrh2a4;
	wire			Csh2a4;
	wire			Jsh2a4;
	wire			Qsh2a4;
	wire			Xsh2a4;
	wire			Eth2a4;
	wire			Lth2a4;
	wire			Sth2a4;
	wire			Zth2a4;
	wire			Guh2a4;
	wire			Nuh2a4;
	wire			Uuh2a4;
	wire			Bvh2a4;
	wire			Ivh2a4;
	wire			Pvh2a4;
	wire			Wvh2a4;
	wire			Dwh2a4;
	wire			Kwh2a4;
	wire			Rwh2a4;
	wire			Ywh2a4;
	wire			Fxh2a4;
	wire			Mxh2a4;
	wire			Txh2a4;
	wire			Ayh2a4;
	wire			Hyh2a4;
	wire			Oyh2a4;
	wire			Vyh2a4;
	wire			Czh2a4;
	wire			Jzh2a4;
	wire			Qzh2a4;
	wire			Xzh2a4;
	wire			E0i2a4;
	wire			L0i2a4;
	wire			S0i2a4;
	wire			Z0i2a4;
	wire			G1i2a4;
	wire			N1i2a4;
	wire			U1i2a4;
	wire			B2i2a4;
	wire			I2i2a4;
	wire			P2i2a4;
	wire			W2i2a4;
	wire			D3i2a4;
	wire			K3i2a4;
	wire			R3i2a4;
	wire			Y3i2a4;
	wire			F4i2a4;
	wire			M4i2a4;
	wire			T4i2a4;
	wire			A5i2a4;
	wire			H5i2a4;
	wire			O5i2a4;
	wire			V5i2a4;
	wire			C6i2a4;
	wire			J6i2a4;
	wire			Q6i2a4;
	wire			X6i2a4;
	wire			E7i2a4;
	wire			L7i2a4;
	wire			S7i2a4;
	wire			Z7i2a4;
	wire			G8i2a4;
	wire			N8i2a4;
	wire			U8i2a4;
	wire			B9i2a4;
	wire			I9i2a4;
	wire			P9i2a4;
	wire			W9i2a4;
	wire			Dai2a4;
	wire			Kai2a4;
	wire			Rai2a4;
	wire			Yai2a4;
	wire			Fbi2a4;
	wire			Mbi2a4;
	wire			Tbi2a4;
	wire			Aci2a4;
	wire			Hci2a4;
	wire			Oci2a4;
	wire			Vci2a4;
	wire			Cdi2a4;
	wire			Jdi2a4;
	wire			Qdi2a4;
	wire			Xdi2a4;
	wire			Eei2a4;
	wire			Lei2a4;
	wire			Sei2a4;
	wire			Zei2a4;
	wire			Gfi2a4;
	wire			Nfi2a4;
	wire			Ufi2a4;
	wire			Bgi2a4;
	wire			Igi2a4;
	wire			Pgi2a4;
	wire			Wgi2a4;
	wire			Dhi2a4;
	wire			Khi2a4;
	wire			Rhi2a4;
	wire			Yhi2a4;
	wire			Fii2a4;
	wire			Mii2a4;
	wire			Tii2a4;
	wire			Aji2a4;
	wire			Hji2a4;
	wire			Oji2a4;
	wire			Vji2a4;
	wire			Cki2a4;
	wire			Jki2a4;
	wire			Qki2a4;
	wire			Xki2a4;
	wire			Eli2a4;
	wire			Lli2a4;
	wire			Sli2a4;
	wire			Zli2a4;
	wire			Gmi2a4;
	wire			Nmi2a4;
	wire			Umi2a4;
	wire			Bni2a4;
	wire			Ini2a4;
	wire			Pni2a4;
	wire			Wni2a4;
	wire			Doi2a4;
	wire			Koi2a4;
	wire			Roi2a4;
	wire			Yoi2a4;
	wire			Fpi2a4;
	wire			Mpi2a4;
	wire			Tpi2a4;
	wire			Aqi2a4;
	wire			Hqi2a4;
	wire			Oqi2a4;
	wire			Vqi2a4;
	wire			Cri2a4;
	wire			Jri2a4;
	wire			Qri2a4;
	wire			Xri2a4;
	wire			Esi2a4;
	wire			Lsi2a4;
	wire			Ssi2a4;
	wire			Zsi2a4;
	wire			Gti2a4;
	wire			Nti2a4;
	wire			Uti2a4;
	wire			Bui2a4;
	wire			Iui2a4;
	wire			Pui2a4;
	wire			Wui2a4;
	wire			Dvi2a4;
	wire			Kvi2a4;
	wire			Rvi2a4;
	wire			Yvi2a4;
	wire			Fwi2a4;
	wire			Mwi2a4;
	wire			Twi2a4;
	wire			Axi2a4;
	wire			Hxi2a4;
	wire			Oxi2a4;
	wire			Vxi2a4;
	wire			Cyi2a4;
	wire			Jyi2a4;
	wire			Qyi2a4;
	wire			Xyi2a4;
	wire			Ezi2a4;
	wire			Lzi2a4;
	wire			Szi2a4;
	wire			Zzi2a4;
	wire			G0j2a4;
	wire			N0j2a4;
	wire			U0j2a4;
	wire			B1j2a4;
	wire			I1j2a4;
	wire			P1j2a4;
	wire			W1j2a4;
	wire			D2j2a4;
	wire			K2j2a4;
	wire			R2j2a4;
	wire			Y2j2a4;
	wire			F3j2a4;
	wire			M3j2a4;
	wire			T3j2a4;
	wire			A4j2a4;
	wire			H4j2a4;
	wire			O4j2a4;
	wire			V4j2a4;
	wire			C5j2a4;
	wire			J5j2a4;
	wire			Q5j2a4;
	wire			X5j2a4;
	wire			E6j2a4;
	wire			L6j2a4;
	wire			S6j2a4;
	wire			Z6j2a4;
	wire			G7j2a4;
	wire			N7j2a4;
	wire			U7j2a4;
	wire			B8j2a4;
	wire			I8j2a4;
	wire			P8j2a4;
	wire			W8j2a4;
	wire			D9j2a4;
	wire			K9j2a4;
	wire			R9j2a4;
	wire			Y9j2a4;
	wire			Faj2a4;
	wire			Maj2a4;
	wire			Taj2a4;
	wire			Abj2a4;
	wire			Hbj2a4;
	wire			Obj2a4;
	wire			Vbj2a4;
	wire			Ccj2a4;
	wire			Jcj2a4;
	wire			Qcj2a4;
	wire			Xcj2a4;
	wire			Edj2a4;
	wire			Ldj2a4;
	wire			Sdj2a4;
	wire			Zdj2a4;
	wire			Gej2a4;
	wire			Nej2a4;
	wire			Uej2a4;
	wire			Bfj2a4;
	wire			Ifj2a4;
	wire			Pfj2a4;
	wire			Wfj2a4;
	wire			Dgj2a4;
	wire			Kgj2a4;
	wire			Rgj2a4;
	wire			Ygj2a4;
	wire			Fhj2a4;
	wire			Mhj2a4;
	wire			Thj2a4;
	wire			Aij2a4;
	wire			Hij2a4;
	wire			Oij2a4;
	wire			Vij2a4;
	wire			Cjj2a4;
	wire			Jjj2a4;
	wire			Qjj2a4;
	wire			Xjj2a4;
	wire			Ekj2a4;
	wire			Lkj2a4;
	wire			Skj2a4;
	wire			Zkj2a4;
	wire			Glj2a4;
	wire			Nlj2a4;
	wire			Ulj2a4;
	wire			Bmj2a4;
	wire			Imj2a4;
	wire			Pmj2a4;
	wire			Wmj2a4;
	wire			Dnj2a4;
	wire			Knj2a4;
	wire			Rnj2a4;
	wire			Ynj2a4;
	wire			Foj2a4;
	wire			Moj2a4;
	wire			Toj2a4;
	wire			Apj2a4;
	wire			Hpj2a4;
	wire			Opj2a4;
	wire			Vpj2a4;
	wire			Cqj2a4;
	wire			Jqj2a4;
	wire			Qqj2a4;
	wire			Xqj2a4;
	wire			Erj2a4;
	wire			Lrj2a4;
	wire			Srj2a4;
	wire			Zrj2a4;
	wire			Gsj2a4;
	wire			Nsj2a4;
	wire			Usj2a4;
	wire			Btj2a4;
	wire			Itj2a4;
	wire			Ptj2a4;
	wire			Wtj2a4;
	wire			Duj2a4;
	wire			Kuj2a4;
	wire			Ruj2a4;
	wire			Yuj2a4;
	wire			Fvj2a4;
	wire			Mvj2a4;
	wire			Tvj2a4;
	wire			Awj2a4;
	wire			Hwj2a4;
	wire			Owj2a4;
	wire			Vwj2a4;
	wire			Cxj2a4;
	wire			Jxj2a4;
	wire			Qxj2a4;
	wire			Xxj2a4;
	wire			Eyj2a4;
	wire			Lyj2a4;
	wire			Syj2a4;
	wire			Zyj2a4;
	wire			Gzj2a4;
	wire			Nzj2a4;
	wire			Uzj2a4;
	wire			B0k2a4;
	wire			I0k2a4;
	wire			P0k2a4;
	wire			W0k2a4;
	wire			D1k2a4;
	wire			K1k2a4;
	wire			R1k2a4;
	wire			Y1k2a4;
	wire			F2k2a4;
	wire			M2k2a4;
	wire			T2k2a4;
	wire			A3k2a4;
	wire			H3k2a4;
	wire			O3k2a4;
	wire			V3k2a4;
	wire			C4k2a4;
	wire			J4k2a4;
	wire			Q4k2a4;
	wire			X4k2a4;
	wire			E5k2a4;
	wire			L5k2a4;
	wire			S5k2a4;
	wire			Z5k2a4;
	wire			G6k2a4;
	wire			N6k2a4;
	wire			U6k2a4;
	wire			B7k2a4;
	wire			I7k2a4;
	wire			P7k2a4;
	wire			W7k2a4;
	wire			D8k2a4;
	wire			K8k2a4;
	wire			R8k2a4;
	wire			Y8k2a4;
	wire			F9k2a4;
	wire			M9k2a4;
	wire			T9k2a4;
	wire			Aak2a4;
	wire			Hak2a4;
	wire			Oak2a4;
	wire			Vak2a4;
	wire			Cbk2a4;
	wire			Jbk2a4;
	wire			Qbk2a4;
	wire			Xbk2a4;
	wire			Eck2a4;
	wire			Lck2a4;
	wire			Sck2a4;
	wire			Zck2a4;
	wire			Gdk2a4;
	wire			Ndk2a4;
	wire			Udk2a4;
	wire			Bek2a4;
	wire			Iek2a4;
	wire			Pek2a4;
	wire			Wek2a4;
	wire			Dfk2a4;
	wire			Kfk2a4;
	wire			Rfk2a4;
	wire			Yfk2a4;
	wire			Fgk2a4;
	wire			Mgk2a4;
	wire			Tgk2a4;
	wire			Ahk2a4;
	wire			Hhk2a4;
	wire			Ohk2a4;
	wire			Vhk2a4;
	wire			Cik2a4;
	wire			Jik2a4;
	wire			Qik2a4;
	wire			Xik2a4;
	wire			Ejk2a4;
	wire			Ljk2a4;
	wire			Sjk2a4;
	wire			Zjk2a4;
	wire			Gkk2a4;
	wire			Nkk2a4;
	wire			Ukk2a4;
	wire			Blk2a4;
	wire			Ilk2a4;
	wire			Plk2a4;
	wire			Wlk2a4;
	wire			Dmk2a4;
	wire			Kmk2a4;
	wire			Rmk2a4;
	wire			Ymk2a4;
	wire			Fnk2a4;
	wire			Mnk2a4;
	wire			Tnk2a4;
	wire			Aok2a4;
	wire			Hok2a4;
	wire			Ook2a4;
	wire			Vok2a4;
	wire			Cpk2a4;
	wire			Jpk2a4;
	wire			Qpk2a4;
	wire			Xpk2a4;
	wire			Eqk2a4;
	wire			Lqk2a4;
	wire			Sqk2a4;
	wire			Zqk2a4;
	wire			Grk2a4;
	wire			Nrk2a4;
	wire			Urk2a4;
	wire			Bsk2a4;
	wire			Isk2a4;
	wire			Psk2a4;
	wire			Wsk2a4;
	wire			Dtk2a4;
	wire			Ktk2a4;
	wire			Rtk2a4;
	wire			Ytk2a4;
	wire			Fuk2a4;
	wire			Muk2a4;
	wire			Tuk2a4;
	wire			Avk2a4;
	wire			Hvk2a4;
	wire			Ovk2a4;
	wire			Vvk2a4;
	wire			Cwk2a4;
	wire			Jwk2a4;
	wire			Qwk2a4;
	wire			Xwk2a4;
	wire			Exk2a4;
	wire			Lxk2a4;
	wire			Sxk2a4;
	wire			Zxk2a4;
	wire			Gyk2a4;
	wire			Nyk2a4;
	wire			Uyk2a4;
	wire			Bzk2a4;
	wire			Izk2a4;
	wire			Pzk2a4;
	wire			Wzk2a4;
	wire			D0l2a4;
	wire			K0l2a4;
	wire			R0l2a4;
	wire			Y0l2a4;
	wire			F1l2a4;
	wire			M1l2a4;
	wire			T1l2a4;
	wire			A2l2a4;
	wire			H2l2a4;
	wire			O2l2a4;
	wire			V2l2a4;
	wire			C3l2a4;
	wire			J3l2a4;
	wire			Q3l2a4;
	wire			X3l2a4;
	wire			E4l2a4;
	wire			L4l2a4;
	wire			S4l2a4;
	wire			Z4l2a4;
	wire			G5l2a4;
	wire			N5l2a4;
	wire			U5l2a4;
	wire			B6l2a4;
	wire			I6l2a4;
	wire			P6l2a4;
	wire			W6l2a4;
	wire			D7l2a4;
	wire			K7l2a4;
	wire			R7l2a4;
	wire			Y7l2a4;
	wire			F8l2a4;
	wire			M8l2a4;
	wire			T8l2a4;
	wire			A9l2a4;
	wire			H9l2a4;
	wire			O9l2a4;
	wire			V9l2a4;
	wire			Cal2a4;
	wire			Jal2a4;
	wire			Qal2a4;
	wire			Xal2a4;
	wire			Ebl2a4;
	wire			Lbl2a4;
	wire			Sbl2a4;
	wire			Zbl2a4;
	wire			Gcl2a4;
	wire			Ncl2a4;
	wire			Ucl2a4;
	wire			Bdl2a4;
	wire			Idl2a4;
	wire			Pdl2a4;
	wire			Wdl2a4;
	wire			Del2a4;
	wire			Kel2a4;
	wire			Rel2a4;
	wire			Yel2a4;
	wire			Ffl2a4;
	wire			Mfl2a4;
	wire			Tfl2a4;
	wire			Agl2a4;
	wire			Hgl2a4;
	wire			Ogl2a4;
	wire			Vgl2a4;
	wire			Chl2a4;
	wire			Jhl2a4;
	wire			Qhl2a4;
	wire			Xhl2a4;
	wire			Eil2a4;
	wire			Lil2a4;
	wire			Sil2a4;
	wire			Zil2a4;
	wire			Gjl2a4;
	wire			Njl2a4;
	wire			Ujl2a4;
	wire			Bkl2a4;
	wire			Ikl2a4;
	wire			Pkl2a4;
	wire			Wkl2a4;
	wire			Dll2a4;
	wire			Kll2a4;
	wire			Rll2a4;
	wire			Yll2a4;
	wire			Fml2a4;
	wire			Mml2a4;
	wire			Tml2a4;
	wire			Anl2a4;
	wire			Hnl2a4;
	wire			Onl2a4;
	wire			Vnl2a4;
	wire			Col2a4;
	wire			Jol2a4;
	wire			Qol2a4;
	wire			Xol2a4;
	wire			Epl2a4;
	wire			Lpl2a4;
	wire			Spl2a4;
	wire			Zpl2a4;
	wire			Gql2a4;
	wire			Nql2a4;
	wire			Uql2a4;
	wire			Brl2a4;
	wire			Irl2a4;
	wire			Prl2a4;
	wire			Wrl2a4;
	wire			Dsl2a4;
	wire			Ksl2a4;
	wire			Rsl2a4;
	wire			Ysl2a4;
	wire			Ftl2a4;
	wire			Mtl2a4;
	wire			Ttl2a4;
	wire			Aul2a4;
	wire			Hul2a4;
	wire			Oul2a4;
	wire			Vul2a4;
	wire			Cvl2a4;
	wire			Jvl2a4;
	wire			Qvl2a4;
	wire			Xvl2a4;
	wire			Ewl2a4;
	wire			Lwl2a4;
	wire			Swl2a4;
	wire			Zwl2a4;
	wire			Gxl2a4;
	wire			Nxl2a4;
	wire			Uxl2a4;
	wire			Byl2a4;
	wire			Iyl2a4;
	wire			Pyl2a4;
	wire			Wyl2a4;
	wire			Dzl2a4;
	wire			Kzl2a4;
	wire			Rzl2a4;
	wire			Yzl2a4;
	wire			F0m2a4;
	wire			M0m2a4;
	wire			T0m2a4;
	wire			A1m2a4;
	wire			H1m2a4;
	wire			O1m2a4;
	wire			V1m2a4;
	wire			C2m2a4;
	wire			J2m2a4;
	wire			Q2m2a4;
	wire			X2m2a4;
	wire			E3m2a4;
	wire			L3m2a4;
	wire			S3m2a4;
	wire			Z3m2a4;
	wire			G4m2a4;
	wire			N4m2a4;
	wire			U4m2a4;
	wire			B5m2a4;
	wire			I5m2a4;
	wire			P5m2a4;
	wire			W5m2a4;
	wire			D6m2a4;
	wire			K6m2a4;
	wire			R6m2a4;
	wire			Y6m2a4;
	wire			F7m2a4;
	wire			M7m2a4;
	wire			T7m2a4;
	wire			A8m2a4;
	wire			H8m2a4;
	wire			O8m2a4;
	wire			V8m2a4;
	wire			C9m2a4;
	wire			J9m2a4;
	wire			Q9m2a4;
	wire			X9m2a4;
	wire			Eam2a4;
	wire			Lam2a4;
	wire			Sam2a4;
	wire			Zam2a4;
	wire			Gbm2a4;
	wire			Nbm2a4;
	wire			Ubm2a4;
	wire			Bcm2a4;
	wire			Icm2a4;
	wire			Pcm2a4;
	wire			Wcm2a4;
	wire			Ddm2a4;
	wire			Kdm2a4;
	wire			Rdm2a4;
	wire			Ydm2a4;
	wire			Fem2a4;
	wire			Mem2a4;
	wire			Tem2a4;
	wire			Afm2a4;
	wire			Hfm2a4;
	wire			Ofm2a4;
	wire			Vfm2a4;
	wire			Cgm2a4;
	wire			Jgm2a4;
	wire			Qgm2a4;
	wire			Xgm2a4;
	wire			Ehm2a4;
	wire			Lhm2a4;
	wire			Shm2a4;
	wire			Zhm2a4;
	wire			Gim2a4;
	wire			Nim2a4;
	wire			Uim2a4;
	wire			Bjm2a4;
	wire			Ijm2a4;
	wire			Pjm2a4;
	wire			Wjm2a4;
	wire			Dkm2a4;
	wire			Kkm2a4;
	wire			Rkm2a4;
	wire			Ykm2a4;
	wire			Flm2a4;
	wire			Mlm2a4;
	wire			Tlm2a4;
	wire			Amm2a4;
	wire			Hmm2a4;
	wire			Omm2a4;
	wire			Vmm2a4;
	wire			Cnm2a4;
	wire			Jnm2a4;
	wire			Qnm2a4;
	wire			Xnm2a4;
	wire			Eom2a4;
	wire			Lom2a4;
	wire			Som2a4;
	wire			Zom2a4;
	wire			Gpm2a4;
	wire			Npm2a4;
	wire			Upm2a4;
	wire			Bqm2a4;
	wire			Iqm2a4;
	wire			Pqm2a4;
	wire			Wqm2a4;
	wire			Drm2a4;
	wire			Krm2a4;
	wire			Rrm2a4;
	wire			Yrm2a4;
	wire			Fsm2a4;
	wire			Msm2a4;
	wire			Tsm2a4;
	wire			Atm2a4;
	wire			Htm2a4;
	wire			Otm2a4;
	wire			Vtm2a4;
	wire			Cum2a4;
	wire			Jum2a4;
	wire			Qum2a4;
	wire			Xum2a4;
	wire			Evm2a4;
	wire			Lvm2a4;
	wire			Svm2a4;
	wire			Zvm2a4;
	wire			Gwm2a4;
	wire			Nwm2a4;
	wire			Uwm2a4;
	wire			Bxm2a4;
	wire			Ixm2a4;
	wire			Pxm2a4;
	wire			Wxm2a4;
	wire			Dym2a4;
	wire			Kym2a4;
	wire			Rym2a4;
	wire			Yym2a4;
	wire			Fzm2a4;
	wire			Mzm2a4;
	wire			Tzm2a4;
	wire			A0n2a4;
	wire			H0n2a4;
	wire			O0n2a4;
	wire			V0n2a4;
	wire			C1n2a4;
	wire			J1n2a4;
	wire			Q1n2a4;
	wire			X1n2a4;
	wire			E2n2a4;
	wire			L2n2a4;
	wire			S2n2a4;
	wire			Z2n2a4;
	wire			G3n2a4;
	wire			N3n2a4;
	wire			U3n2a4;
	wire			B4n2a4;
	wire			I4n2a4;
	wire			P4n2a4;
	wire			W4n2a4;
	wire			D5n2a4;
	wire			K5n2a4;
	wire			R5n2a4;
	wire			Y5n2a4;
	wire			F6n2a4;
	wire			M6n2a4;
	wire			T6n2a4;
	wire			A7n2a4;
	wire			H7n2a4;
	wire			O7n2a4;
	wire			V7n2a4;
	wire			C8n2a4;
	wire			J8n2a4;
	wire			Q8n2a4;
	wire			X8n2a4;
	wire			E9n2a4;
	wire			L9n2a4;
	wire			S9n2a4;
	wire			Z9n2a4;
	wire			Gan2a4;
	wire			Nan2a4;
	wire			Uan2a4;
	wire			Bbn2a4;
	wire			Ibn2a4;
	wire			Pbn2a4;
	wire			Wbn2a4;
	wire			Dcn2a4;
	wire			Kcn2a4;
	wire			Rcn2a4;
	wire			Ycn2a4;
	wire			Fdn2a4;
	wire			Mdn2a4;
	wire			Tdn2a4;
	wire			Aen2a4;
	wire			Hen2a4;
	wire			Oen2a4;
	wire			Ven2a4;
	wire			Cfn2a4;
	wire			Jfn2a4;
	wire			Qfn2a4;
	wire			Xfn2a4;
	wire			Egn2a4;
	wire			Lgn2a4;
	wire			Sgn2a4;
	wire			Zgn2a4;
	wire			Ghn2a4;
	wire			Nhn2a4;
	wire			Uhn2a4;
	wire			Bin2a4;
	wire			Iin2a4;
	wire			Pin2a4;
	wire			Win2a4;
	wire			Djn2a4;
	wire			Kjn2a4;
	wire			Rjn2a4;
	wire			Yjn2a4;
	wire			Fkn2a4;
	wire			Mkn2a4;
	wire			Tkn2a4;
	wire			Aln2a4;
	wire			Hln2a4;
	wire			Oln2a4;
	wire			Vln2a4;
	wire			Cmn2a4;
	wire			Jmn2a4;
	wire			Qmn2a4;
	wire			Xmn2a4;
	wire			Enn2a4;
	wire			Lnn2a4;
	wire			Snn2a4;
	wire			Znn2a4;
	wire			Gon2a4;
	wire			Non2a4;
	wire			Uon2a4;
	wire			Bpn2a4;
	wire			Ipn2a4;
	wire			Ppn2a4;
	wire			Wpn2a4;
	wire			Dqn2a4;
	wire			Kqn2a4;
	wire			Rqn2a4;
	wire			Yqn2a4;
	wire			Frn2a4;
	wire			Mrn2a4;
	wire			Trn2a4;
	wire			Asn2a4;
	wire			Hsn2a4;
	wire			Osn2a4;
	wire			Vsn2a4;
	wire			Ctn2a4;
	wire			Jtn2a4;
	wire			Qtn2a4;
	wire			Xtn2a4;
	wire			Eun2a4;
	wire			Lun2a4;
	wire			Sun2a4;
	wire			Zun2a4;
	wire			Gvn2a4;
	wire			Nvn2a4;
	wire			Uvn2a4;
	wire			Bwn2a4;
	wire			Iwn2a4;
	wire			Pwn2a4;
	wire			Wwn2a4;
	wire			Dxn2a4;
	wire			Kxn2a4;
	wire			Rxn2a4;
	wire			Yxn2a4;
	wire			Fyn2a4;
	wire			Myn2a4;
	wire			Tyn2a4;
	wire			Azn2a4;
	wire			Hzn2a4;
	wire			Ozn2a4;
	wire			Vzn2a4;
	wire			C0o2a4;
	wire			J0o2a4;
	wire			Q0o2a4;
	wire			X0o2a4;
	wire			E1o2a4;
	wire			L1o2a4;
	wire			S1o2a4;
	wire			Z1o2a4;
	wire			G2o2a4;
	wire			N2o2a4;
	wire			U2o2a4;
	wire			B3o2a4;
	wire			I3o2a4;
	wire			P3o2a4;
	wire			W3o2a4;
	wire			D4o2a4;
	wire			K4o2a4;
	wire			R4o2a4;
	wire			Y4o2a4;
	wire			F5o2a4;
	wire			M5o2a4;
	wire			T5o2a4;
	wire			A6o2a4;
	wire			H6o2a4;
	wire			O6o2a4;
	wire			V6o2a4;
	wire			C7o2a4;
	wire			J7o2a4;
	wire			Q7o2a4;
	wire			X7o2a4;
	wire			E8o2a4;
	wire			L8o2a4;
	wire			S8o2a4;
	wire			Z8o2a4;
	wire			G9o2a4;
	wire			N9o2a4;
	wire			U9o2a4;
	wire			Bao2a4;
	wire			Iao2a4;
	wire			Pao2a4;
	wire			Wao2a4;
	wire			Dbo2a4;
	wire			Kbo2a4;
	wire			Rbo2a4;
	wire			Ybo2a4;
	wire			Fco2a4;
	wire			Mco2a4;
	wire			Tco2a4;
	wire			Ado2a4;
	wire			Hdo2a4;
	wire			Odo2a4;
	wire			Vdo2a4;
	wire			Ceo2a4;
	wire			Jeo2a4;
	wire			Qeo2a4;
	wire			Xeo2a4;
	wire			Efo2a4;
	wire			Lfo2a4;
	wire			Sfo2a4;
	wire			Zfo2a4;
	wire			Ggo2a4;
	wire			Ngo2a4;
	wire			Ugo2a4;
	wire			Bho2a4;
	wire			Iho2a4;
	wire			Pho2a4;
	wire			Who2a4;
	wire			Dio2a4;
	wire			Kio2a4;
	wire			Rio2a4;
	wire			Yio2a4;
	wire			Fjo2a4;
	wire			Mjo2a4;
	wire			Tjo2a4;
	wire			Ako2a4;
	wire			Hko2a4;
	wire			Oko2a4;
	wire			Vko2a4;
	wire			Clo2a4;
	wire			Jlo2a4;
	wire			Qlo2a4;
	wire			Xlo2a4;
	wire			Emo2a4;
	wire			Lmo2a4;
	wire			Smo2a4;
	wire			Zmo2a4;
	wire			Gno2a4;
	wire			Nno2a4;
	wire			Uno2a4;
	wire			Boo2a4;
	wire			Ioo2a4;
	wire			Poo2a4;
	wire			Woo2a4;
	wire			Dpo2a4;
	wire			Kpo2a4;
	wire			Rpo2a4;
	wire			Ypo2a4;
	wire			Fqo2a4;
	wire			Mqo2a4;
	wire			Tqo2a4;
	wire			Aro2a4;
	wire			Hro2a4;
	wire			Oro2a4;
	wire			Vro2a4;
	wire			Cso2a4;
	wire			Jso2a4;
	wire			Qso2a4;
	wire			Xso2a4;
	wire			Eto2a4;
	wire			Lto2a4;
	wire			Sto2a4;
	wire			Zto2a4;
	wire			Guo2a4;
	wire			Nuo2a4;
	wire			Uuo2a4;
	wire			Bvo2a4;
	wire			Ivo2a4;
	wire			Pvo2a4;
	wire			Wvo2a4;
	wire			Dwo2a4;
	wire			Kwo2a4;
	wire			Rwo2a4;
	wire			Ywo2a4;
	wire			Fxo2a4;
	wire			Mxo2a4;
	wire			Txo2a4;
	wire			Ayo2a4;
	wire			Hyo2a4;
	wire			Oyo2a4;
	wire			Vyo2a4;
	wire			Czo2a4;
	wire			Jzo2a4;
	wire			Qzo2a4;
	wire			Xzo2a4;
	wire			E0p2a4;
	wire			L0p2a4;
	wire			S0p2a4;
	wire			Z0p2a4;
	wire			G1p2a4;
	wire			N1p2a4;
	wire			U1p2a4;
	wire			B2p2a4;
	wire			I2p2a4;
	wire			P2p2a4;
	wire			W2p2a4;
	wire			D3p2a4;
	wire			K3p2a4;
	wire			R3p2a4;
	wire			Y3p2a4;
	wire			F4p2a4;
	wire			M4p2a4;
	wire			T4p2a4;
	wire			A5p2a4;
	wire			H5p2a4;
	wire			O5p2a4;
	wire			V5p2a4;
	wire			C6p2a4;
	wire			J6p2a4;
	wire			Q6p2a4;
	wire			X6p2a4;
	wire			E7p2a4;
	wire			L7p2a4;
	wire			S7p2a4;
	wire			Z7p2a4;
	wire			G8p2a4;
	wire			N8p2a4;
	wire			U8p2a4;
	wire			B9p2a4;
	wire			I9p2a4;
	wire			P9p2a4;
	wire			W9p2a4;
	wire			Dap2a4;
	wire			Kap2a4;
	wire			Rap2a4;
	wire			Yap2a4;
	wire			Fbp2a4;
	wire			Mbp2a4;
	wire			Tbp2a4;
	wire			Acp2a4;
	wire			Hcp2a4;
	wire			Ocp2a4;
	wire			Vcp2a4;
	wire			Cdp2a4;
	wire			Jdp2a4;
	wire			Qdp2a4;
	wire			Xdp2a4;
	wire			Eep2a4;
	wire			Lep2a4;
	wire			Sep2a4;
	wire			Zep2a4;
	wire			Gfp2a4;
	wire			Nfp2a4;
	wire			Ufp2a4;
	wire			Bgp2a4;
	wire			Igp2a4;
	wire			Pgp2a4;
	wire			Wgp2a4;
	wire			Dhp2a4;
	wire			Khp2a4;
	wire			Rhp2a4;
	wire			Yhp2a4;
	wire			Fip2a4;
	wire			Mip2a4;
	wire			Tip2a4;
	wire			Ajp2a4;
	wire			Hjp2a4;
	wire			Ojp2a4;
	wire			Vjp2a4;
	wire			Ckp2a4;
	wire			Jkp2a4;
	wire			Qkp2a4;
	wire			Xkp2a4;
	wire			Elp2a4;
	wire			Llp2a4;
	wire			Slp2a4;
	wire			Zlp2a4;
	wire			Gmp2a4;
	wire			Nmp2a4;
	wire			Ump2a4;
	wire			Bnp2a4;
	wire			Inp2a4;
	wire			Pnp2a4;
	wire			Wnp2a4;
	wire			Dop2a4;
	wire			Kop2a4;
	wire			Rop2a4;
	wire			Yop2a4;
	wire			Fpp2a4;
	wire			Mpp2a4;
	wire			Tpp2a4;
	wire			Aqp2a4;
	wire			Hqp2a4;
	wire			Oqp2a4;
	wire			Vqp2a4;
	wire			Crp2a4;
	wire			Jrp2a4;
	wire			Qrp2a4;
	wire			Xrp2a4;
	wire			Esp2a4;
	wire			Lsp2a4;
	wire			Ssp2a4;
	wire			Zsp2a4;
	wire			Gtp2a4;
	wire			Ntp2a4;
	wire			Utp2a4;
	wire			Bup2a4;
	wire			Iup2a4;
	wire			Pup2a4;
	wire			Wup2a4;
	wire			Dvp2a4;
	wire			Kvp2a4;
	wire			Rvp2a4;
	wire			Yvp2a4;
	wire			Fwp2a4;
	wire			Mwp2a4;
	wire			Twp2a4;
	wire			Axp2a4;
	wire			Hxp2a4;
	wire			Oxp2a4;
	wire			Vxp2a4;
	wire			Cyp2a4;
	wire			Jyp2a4;
	wire			Qyp2a4;
	wire			Xyp2a4;
	wire			Ezp2a4;
	wire			Lzp2a4;
	wire			Szp2a4;
	wire			Zzp2a4;
	wire			G0q2a4;
	wire			N0q2a4;
	wire			U0q2a4;
	wire			B1q2a4;
	wire			I1q2a4;
	wire			P1q2a4;
	wire			W1q2a4;
	wire			D2q2a4;
	wire			K2q2a4;
	wire			R2q2a4;
	wire			Y2q2a4;
	wire			F3q2a4;
	wire			M3q2a4;
	wire			T3q2a4;
	wire			A4q2a4;
	wire			H4q2a4;
	wire			O4q2a4;
	wire			V4q2a4;
	wire			C5q2a4;
	wire			J5q2a4;
	wire			Q5q2a4;
	wire			X5q2a4;
	wire			E6q2a4;
	wire			L6q2a4;
	wire			S6q2a4;
	wire			Z6q2a4;
	wire			G7q2a4;
	wire			N7q2a4;
	wire			U7q2a4;
	wire			B8q2a4;
	wire			I8q2a4;
	wire			P8q2a4;
	wire			W8q2a4;
	wire			D9q2a4;
	wire			K9q2a4;
	wire			R9q2a4;
	wire			Y9q2a4;
	wire			Faq2a4;
	wire			Maq2a4;
	wire			Taq2a4;
	wire			Abq2a4;
	wire			Hbq2a4;
	wire			Obq2a4;
	wire			Vbq2a4;
	wire			Ccq2a4;
	wire			Jcq2a4;
	wire			Qcq2a4;
	wire			Xcq2a4;
	wire			Edq2a4;
	wire			Ldq2a4;
	wire			Sdq2a4;
	wire			Zdq2a4;
	wire			Geq2a4;
	wire			Neq2a4;
	wire			Ueq2a4;
	wire			Bfq2a4;
	wire			Ifq2a4;
	wire			Pfq2a4;
	wire			Wfq2a4;
	wire			Dgq2a4;
	wire			Kgq2a4;
	wire			Rgq2a4;
	wire			Ygq2a4;
	wire			Fhq2a4;
	wire			Mhq2a4;
	wire			Thq2a4;
	wire			Aiq2a4;
	wire			Hiq2a4;
	wire			Oiq2a4;
	wire			Viq2a4;
	wire			Cjq2a4;
	wire			Jjq2a4;
	wire			Qjq2a4;
	wire			Xjq2a4;
	wire			Ekq2a4;
	wire			Lkq2a4;
	wire			Skq2a4;
	wire			Zkq2a4;
	wire			Glq2a4;
	wire			Nlq2a4;
	wire			Ulq2a4;
	wire			Bmq2a4;
	wire			Imq2a4;
	wire			Pmq2a4;
	wire			Wmq2a4;
	wire			Dnq2a4;
	wire			Knq2a4;
	wire			Rnq2a4;
	wire			Ynq2a4;
	wire			Foq2a4;
	wire			Moq2a4;
	wire			Toq2a4;
	wire			Apq2a4;
	wire			Hpq2a4;
	wire			Opq2a4;
	wire			Vpq2a4;
	wire			Cqq2a4;
	wire			Jqq2a4;
	wire			Qqq2a4;
	wire			Xqq2a4;
	wire			Erq2a4;
	wire			Lrq2a4;
	wire			Srq2a4;
	wire			Zrq2a4;
	wire			Gsq2a4;
	wire			Nsq2a4;
	wire			Usq2a4;
	wire			Btq2a4;
	wire			Itq2a4;
	wire			Ptq2a4;
	wire			Wtq2a4;
	wire			Duq2a4;
	wire			Kuq2a4;
	wire			Ruq2a4;
	wire			Yuq2a4;
	wire			Fvq2a4;
	wire			Mvq2a4;
	wire			Tvq2a4;
	wire			Awq2a4;
	wire			Hwq2a4;
	wire			Owq2a4;
	wire			Vwq2a4;
	wire			Cxq2a4;
	wire			Jxq2a4;
	wire			Qxq2a4;
	wire			Xxq2a4;
	wire			Eyq2a4;
	wire			Lyq2a4;
	wire			Syq2a4;
	wire			Zyq2a4;
	wire			Gzq2a4;
	wire			Nzq2a4;
	wire			Uzq2a4;
	wire			B0r2a4;
	wire			I0r2a4;
	wire			P0r2a4;
	wire			W0r2a4;
	wire			D1r2a4;
	wire			K1r2a4;
	wire			R1r2a4;
	wire			Y1r2a4;
	wire			F2r2a4;
	wire			M2r2a4;
	wire			T2r2a4;
	wire			A3r2a4;
	wire			H3r2a4;
	wire			O3r2a4;
	wire			V3r2a4;
	wire			C4r2a4;
	wire			J4r2a4;
	wire			Q4r2a4;
	wire			X4r2a4;
	wire			E5r2a4;
	wire			L5r2a4;
	wire			S5r2a4;
	wire			Z5r2a4;
	wire			G6r2a4;
	wire			N6r2a4;
	wire			U6r2a4;
	wire			B7r2a4;
	wire			I7r2a4;
	wire			P7r2a4;
	wire			W7r2a4;
	wire			D8r2a4;
	wire			K8r2a4;
	wire			R8r2a4;
	wire			Y8r2a4;
	wire			F9r2a4;
	wire			M9r2a4;
	wire			T9r2a4;
	wire			Aar2a4;
	wire			Har2a4;
	wire			Oar2a4;
	wire			Var2a4;
	wire			Cbr2a4;
	wire			Jbr2a4;
	wire			Qbr2a4;
	wire			Xbr2a4;
	wire			Ecr2a4;
	wire			Lcr2a4;
	wire			Scr2a4;
	wire			Zcr2a4;
	wire			Gdr2a4;
	wire			Ndr2a4;
	wire			Udr2a4;
	wire			Ber2a4;
	wire			Ier2a4;
	wire			Per2a4;
	wire			Wer2a4;
	wire			Dfr2a4;
	wire			Kfr2a4;
	wire			Rfr2a4;
	wire			Yfr2a4;
	wire			Fgr2a4;
	wire			Mgr2a4;
	wire			Tgr2a4;
	wire			Ahr2a4;
	wire			Hhr2a4;
	wire			Ohr2a4;
	wire			Vhr2a4;
	wire			Cir2a4;
	wire			Jir2a4;
	wire			Qir2a4;
	wire			Xir2a4;
	wire			Ejr2a4;
	wire			Ljr2a4;
	wire			Sjr2a4;
	wire			Zjr2a4;
	wire			Gkr2a4;
	wire			Nkr2a4;
	wire			Ukr2a4;
	wire			Blr2a4;
	wire			Ilr2a4;
	wire			Plr2a4;
	wire			Wlr2a4;
	wire			Dmr2a4;
	wire			Kmr2a4;
	wire			Rmr2a4;
	wire			Ymr2a4;
	wire			Fnr2a4;
	wire			Mnr2a4;
	wire			Tnr2a4;
	wire			Aor2a4;
	wire			Hor2a4;
	wire			Oor2a4;
	wire			Vor2a4;
	wire			Cpr2a4;
	wire			Jpr2a4;
	wire			Qpr2a4;
	wire			Xpr2a4;
	wire			Eqr2a4;
	wire			Lqr2a4;
	wire			Sqr2a4;
	wire			Zqr2a4;
	wire			Grr2a4;
	wire			Nrr2a4;
	wire			Urr2a4;
	wire			Bsr2a4;
	wire			Isr2a4;
	wire			Psr2a4;
	wire			Wsr2a4;
	wire			Dtr2a4;
	wire			Ktr2a4;
	wire			Rtr2a4;
	wire			Ytr2a4;
	wire			Fur2a4;
	wire			Mur2a4;
	wire			Tur2a4;
	wire			Avr2a4;
	wire			Hvr2a4;
	wire			Ovr2a4;
	wire			Vvr2a4;
	wire			Cwr2a4;
	wire			Jwr2a4;
	wire			Qwr2a4;
	wire			Xwr2a4;
	wire			Exr2a4;
	wire			Lxr2a4;
	wire			Sxr2a4;
	wire			Zxr2a4;
	wire			Gyr2a4;
	wire			Nyr2a4;
	wire			Uyr2a4;
	wire			Bzr2a4;
	wire			Izr2a4;
	wire			Pzr2a4;
	wire			Wzr2a4;
	wire			D0s2a4;
	wire			K0s2a4;
	wire			R0s2a4;
	wire			Y0s2a4;
	wire			F1s2a4;
	wire			M1s2a4;
	wire			T1s2a4;
	wire			A2s2a4;
	wire			H2s2a4;
	wire			O2s2a4;
	wire			V2s2a4;
	wire			C3s2a4;
	wire			J3s2a4;
	wire			Q3s2a4;
	wire			X3s2a4;
	wire			E4s2a4;
	wire			L4s2a4;
	wire			S4s2a4;
	wire			Z4s2a4;
	wire			G5s2a4;
	wire			N5s2a4;
	wire			U5s2a4;
	wire			B6s2a4;
	wire			I6s2a4;
	wire			P6s2a4;
	wire			W6s2a4;
	wire			D7s2a4;
	wire			K7s2a4;
	wire			R7s2a4;
	wire			Y7s2a4;
	wire			F8s2a4;
	wire			M8s2a4;
	wire			T8s2a4;
	wire			A9s2a4;
	wire			H9s2a4;
	wire			O9s2a4;
	wire			V9s2a4;
	wire			Cas2a4;
	wire			Jas2a4;
	wire			Qas2a4;
	wire			Xas2a4;
	wire			Ebs2a4;
	wire			Lbs2a4;
	wire			Sbs2a4;
	wire			Zbs2a4;
	wire			Gcs2a4;
	wire			Ncs2a4;
	wire			Ucs2a4;
	wire			Bds2a4;
	wire			Ids2a4;
	wire			Pds2a4;
	wire			Wds2a4;
	wire			Des2a4;
	wire			Kes2a4;
	wire			Res2a4;
	wire			Yes2a4;
	wire			Ffs2a4;
	wire			Mfs2a4;
	wire			Tfs2a4;
	wire			Ags2a4;
	wire			Hgs2a4;
	wire			Ogs2a4;
	wire			Vgs2a4;
	wire			Chs2a4;
	wire			Jhs2a4;
	wire			Qhs2a4;
	wire			Xhs2a4;
	wire			Eis2a4;
	wire			Lis2a4;
	wire			Sis2a4;
	wire			Zis2a4;
	wire			Gjs2a4;
	wire			Njs2a4;
	wire			Ujs2a4;
	wire			Bks2a4;
	wire			Iks2a4;
	wire			Pks2a4;
	wire			Wks2a4;
	wire			Dls2a4;
	wire			Kls2a4;
	wire			Rls2a4;
	wire			Yls2a4;
	wire			Fms2a4;
	wire			Mms2a4;
	wire			Tms2a4;
	wire			Ans2a4;
	wire			Hns2a4;
	wire			Ons2a4;
	wire			Vns2a4;
	wire			Cos2a4;
	wire			Jos2a4;
	wire			Qos2a4;
	wire			Xos2a4;
	wire			Eps2a4;
	wire			Lps2a4;
	wire			Sps2a4;
	wire			Zps2a4;
	wire			Gqs2a4;
	wire			Nqs2a4;
	wire			Uqs2a4;
	wire			Brs2a4;
	wire			Irs2a4;
	wire			Prs2a4;
	wire			Wrs2a4;
	wire			Dss2a4;
	wire			Kss2a4;
	wire			Rss2a4;
	wire			Yss2a4;
	wire			Fts2a4;
	wire			Mts2a4;
	wire			Tts2a4;
	wire			Aus2a4;
	wire			Hus2a4;
	wire			Ous2a4;
	wire			Vus2a4;
	wire			Cvs2a4;
	wire			Jvs2a4;
	wire			Qvs2a4;
	wire			Xvs2a4;
	wire			Ews2a4;
	wire			Lws2a4;
	wire			Sws2a4;
	wire			Zws2a4;
	wire			Gxs2a4;
	wire			Nxs2a4;
	wire			Uxs2a4;
	wire			Bys2a4;
	wire			Iys2a4;
	wire			Pys2a4;
	wire			Wys2a4;
	wire			Dzs2a4;
	wire			Kzs2a4;
	wire			Rzs2a4;
	wire			Yzs2a4;
	wire			F0t2a4;
	wire			M0t2a4;
	wire			T0t2a4;
	wire			A1t2a4;
	wire			H1t2a4;
	wire			O1t2a4;
	wire			V1t2a4;
	wire			C2t2a4;
	wire			J2t2a4;
	wire			Q2t2a4;
	wire			X2t2a4;
	wire			E3t2a4;
	wire			L3t2a4;
	wire			S3t2a4;
	wire			Z3t2a4;
	wire			G4t2a4;
	wire			N4t2a4;
	wire			U4t2a4;
	wire			B5t2a4;
	wire			I5t2a4;
	wire			P5t2a4;
	wire			W5t2a4;
	wire			D6t2a4;
	wire			K6t2a4;
	wire			R6t2a4;
	wire			Y6t2a4;
	wire			F7t2a4;
	wire			M7t2a4;
	wire			T7t2a4;
	wire			A8t2a4;
	wire			H8t2a4;
	wire			O8t2a4;
	wire			V8t2a4;
	wire			C9t2a4;
	wire			J9t2a4;
	wire			Q9t2a4;
	wire			X9t2a4;
	wire			Eat2a4;
	wire			Lat2a4;
	wire			Sat2a4;
	wire			Zat2a4;
	wire			Gbt2a4;
	wire			Nbt2a4;
	wire			Ubt2a4;
	wire			Bct2a4;
	wire			Ict2a4;
	wire			Pct2a4;
	wire			Wct2a4;
	wire			Ddt2a4;
	wire			Kdt2a4;
	wire			Rdt2a4;
	wire			Ydt2a4;
	wire			Fet2a4;
	wire			Met2a4;
	wire			Tet2a4;
	wire			Aft2a4;
	wire			Hft2a4;
	wire			Oft2a4;
	wire			Vft2a4;
	wire			Cgt2a4;
	wire			Jgt2a4;
	wire			Qgt2a4;
	wire			Xgt2a4;
	wire			Eht2a4;
	wire			Lht2a4;
	wire			Sht2a4;
	wire			Zht2a4;
	wire			Git2a4;
	wire			Nit2a4;
	wire			Uit2a4;
	wire			Bjt2a4;
	wire			Ijt2a4;
	wire			Pjt2a4;
	wire			Wjt2a4;
	wire			Dkt2a4;
	wire			Kkt2a4;
	wire			Rkt2a4;
	wire			Ykt2a4;
	wire			Flt2a4;
	wire			Mlt2a4;
	wire			Tlt2a4;
	wire			Amt2a4;
	wire			Hmt2a4;
	wire			Omt2a4;
	wire			Vmt2a4;
	wire			Cnt2a4;
	wire			Jnt2a4;
	wire			Qnt2a4;
	wire			Xnt2a4;
	wire			Eot2a4;
	wire			Lot2a4;
	wire			Sot2a4;
	wire			Zot2a4;
	wire			Gpt2a4;
	wire			Npt2a4;
	wire			Upt2a4;
	wire			Bqt2a4;
	wire			Iqt2a4;
	wire			Pqt2a4;
	wire			Wqt2a4;
	wire			Drt2a4;
	wire			Krt2a4;
	wire			Rrt2a4;
	wire			Yrt2a4;
	wire			Fst2a4;
	wire			Mst2a4;
	wire			Tst2a4;
	wire			Att2a4;
	wire			Htt2a4;
	wire			Ott2a4;
	wire			Vtt2a4;
	wire			Cut2a4;
	wire			Jut2a4;
	wire			Qut2a4;
	wire			Xut2a4;
	wire			Evt2a4;
	wire			Lvt2a4;
	wire			Svt2a4;
	wire			Zvt2a4;
	wire			Gwt2a4;
	wire			Nwt2a4;
	wire			Uwt2a4;
	wire			Bxt2a4;
	wire			Ixt2a4;
	wire			Pxt2a4;
	wire			Wxt2a4;
	wire			Dyt2a4;
	wire			Kyt2a4;
	wire			Ryt2a4;
	wire			Yyt2a4;
	wire			Fzt2a4;
	wire			Mzt2a4;
	wire			Tzt2a4;
	wire			A0u2a4;
	wire			H0u2a4;
	wire			O0u2a4;
	wire			V0u2a4;
	wire			C1u2a4;
	wire			J1u2a4;
	wire			Q1u2a4;
	wire			X1u2a4;
	wire			E2u2a4;
	wire			L2u2a4;
	wire			S2u2a4;
	wire			Z2u2a4;
	wire			G3u2a4;
	wire			N3u2a4;
	wire			U3u2a4;
	wire			B4u2a4;
	wire			I4u2a4;
	wire			P4u2a4;
	wire			W4u2a4;
	wire			D5u2a4;
	wire			K5u2a4;
	wire			R5u2a4;
	wire			Y5u2a4;
	wire			F6u2a4;
	wire			M6u2a4;
	wire			T6u2a4;
	wire			A7u2a4;
	wire			H7u2a4;
	wire			O7u2a4;
	wire			V7u2a4;
	wire			C8u2a4;
	wire			J8u2a4;
	wire			Q8u2a4;
	wire			X8u2a4;
	wire			E9u2a4;
	wire			L9u2a4;
	wire			S9u2a4;
	wire			Z9u2a4;
	wire			Gau2a4;
	wire			Nau2a4;
	wire			Uau2a4;
	wire			Bbu2a4;
	wire			Ibu2a4;
	wire			Pbu2a4;
	wire			Wbu2a4;
	wire			Dcu2a4;
	wire			Kcu2a4;
	wire			Rcu2a4;
	wire			Ycu2a4;
	wire			Fdu2a4;
	wire			Mdu2a4;
	wire			Tdu2a4;
	wire			Aeu2a4;
	wire			Heu2a4;
	wire			Oeu2a4;
	wire			Veu2a4;
	wire			Cfu2a4;
	wire			Jfu2a4;
	wire			Qfu2a4;
	wire			Xfu2a4;
	wire			Egu2a4;
	wire			Lgu2a4;
	wire			Sgu2a4;
	wire			Zgu2a4;
	wire			Ghu2a4;
	wire			Nhu2a4;
	wire			Uhu2a4;
	wire			Biu2a4;
	wire			Iiu2a4;
	wire			Piu2a4;
	wire			Wiu2a4;
	wire			Dju2a4;
	wire			Kju2a4;
	wire			Rju2a4;
	wire			Yju2a4;
	wire			Fku2a4;
	wire			Mku2a4;
	wire			Tku2a4;
	wire			Alu2a4;
	wire			Hlu2a4;
	wire			Olu2a4;
	wire			Vlu2a4;
	wire			Cmu2a4;
	wire			Jmu2a4;
	wire			Qmu2a4;
	wire			Xmu2a4;
	wire			Enu2a4;
	wire			Lnu2a4;
	wire			Snu2a4;
	wire			Znu2a4;
	wire			Gou2a4;
	wire			Nou2a4;
	wire			Uou2a4;
	wire			Bpu2a4;
	wire			Ipu2a4;
	wire			Ppu2a4;
	wire			Wpu2a4;
	wire			Dqu2a4;
	wire			Kqu2a4;
	wire			Rqu2a4;
	wire			Yqu2a4;
	wire			Fru2a4;
	wire			Mru2a4;
	wire			Tru2a4;
	wire			Asu2a4;
	wire			Hsu2a4;
	wire			Osu2a4;
	wire			Vsu2a4;
	wire			Ctu2a4;
	wire			Jtu2a4;
	wire			Qtu2a4;
	wire			Xtu2a4;
	wire			Euu2a4;
	wire			Luu2a4;
	wire			Suu2a4;
	wire			Zuu2a4;
	wire			Gvu2a4;
	wire			Nvu2a4;
	wire			Uvu2a4;
	wire			Bwu2a4;
	wire			Iwu2a4;
	wire			Pwu2a4;
	wire			Wwu2a4;
	wire			Dxu2a4;
	wire			Kxu2a4;
	wire			Rxu2a4;
	wire			Yxu2a4;
	wire			Fyu2a4;
	wire			Myu2a4;
	wire			Tyu2a4;
	wire			Azu2a4;
	wire			Hzu2a4;
	wire			Ozu2a4;
	wire			Vzu2a4;
	wire			C0v2a4;
	wire			J0v2a4;
	wire			Q0v2a4;
	wire			X0v2a4;
	wire			E1v2a4;
	wire			L1v2a4;
	wire			S1v2a4;
	wire			Z1v2a4;
	wire			G2v2a4;
	wire			N2v2a4;
	wire			U2v2a4;
	wire			B3v2a4;
	wire			I3v2a4;
	wire			P3v2a4;
	wire			W3v2a4;
	wire			D4v2a4;
	wire			K4v2a4;
	wire			R4v2a4;
	wire			Y4v2a4;
	wire			F5v2a4;
	wire			M5v2a4;
	wire			T5v2a4;
	wire			A6v2a4;
	wire			H6v2a4;
	wire			O6v2a4;
	wire			V6v2a4;
	wire			C7v2a4;
	wire			J7v2a4;
	wire			Q7v2a4;
	wire			X7v2a4;
	wire			E8v2a4;
	wire			L8v2a4;
	wire			S8v2a4;
	wire			Z8v2a4;
	wire			G9v2a4;
	wire			N9v2a4;
	wire			U9v2a4;
	wire			Bav2a4;
	wire			Iav2a4;
	wire			Pav2a4;
	wire			Wav2a4;
	wire			Dbv2a4;
	wire			Kbv2a4;
	wire			Rbv2a4;
	wire			Ybv2a4;
	wire			Fcv2a4;
	wire			Mcv2a4;
	wire			Tcv2a4;
	wire			Adv2a4;
	wire			Hdv2a4;
	wire			Odv2a4;
	wire			Vdv2a4;
	wire			Cev2a4;
	wire			Jev2a4;
	wire			Qev2a4;
	wire			Xev2a4;
	wire			Efv2a4;
	wire			Lfv2a4;
	wire			Sfv2a4;
	wire			Zfv2a4;
	wire			Ggv2a4;
	wire			Ngv2a4;
	wire			Ugv2a4;
	wire			Bhv2a4;
	wire			Ihv2a4;
	wire			Phv2a4;
	wire			Whv2a4;
	wire			Div2a4;
	wire			Kiv2a4;
	wire			Riv2a4;
	wire			Yiv2a4;
	wire			Fjv2a4;
	wire			Mjv2a4;
	wire			Tjv2a4;
	wire			Akv2a4;
	wire			Hkv2a4;
	wire			Okv2a4;
	wire			Vkv2a4;
	wire			Clv2a4;
	wire			Jlv2a4;
	wire			Qlv2a4;
	wire			Xlv2a4;
	wire			Emv2a4;
	wire			Lmv2a4;
	wire			Smv2a4;
	wire			Zmv2a4;
	wire			Gnv2a4;
	wire			Nnv2a4;
	wire			Unv2a4;
	wire			Bov2a4;
	wire			Iov2a4;
	wire			Pov2a4;
	wire			Wov2a4;
	wire			Dpv2a4;
	wire			Kpv2a4;
	wire			Rpv2a4;
	wire			Ypv2a4;
	wire			Fqv2a4;
	wire			Mqv2a4;
	wire			Tqv2a4;
	wire			Arv2a4;
	wire			Hrv2a4;
	wire			Orv2a4;
	wire			Vrv2a4;
	wire			Csv2a4;
	wire			Jsv2a4;
	wire			Qsv2a4;
	wire			Xsv2a4;
	wire			Etv2a4;
	wire			Ltv2a4;
	wire			Stv2a4;
	wire			Ztv2a4;
	wire			Guv2a4;
	wire			Nuv2a4;
	wire			Uuv2a4;
	wire			Bvv2a4;
	wire			Ivv2a4;
	wire			Pvv2a4;
	wire			Wvv2a4;
	wire			Dwv2a4;
	wire			Kwv2a4;
	wire			Rwv2a4;
	wire			Ywv2a4;
	wire			Fxv2a4;
	wire			Mxv2a4;
	wire			Txv2a4;
	wire			Ayv2a4;
	wire			Hyv2a4;
	wire			Oyv2a4;
	wire			Vyv2a4;
	wire			Czv2a4;
	wire			Jzv2a4;
	wire			Qzv2a4;
	wire			Xzv2a4;
	wire			E0w2a4;
	wire			L0w2a4;
	wire			S0w2a4;
	wire			Z0w2a4;
	wire			G1w2a4;
	wire			N1w2a4;
	wire			U1w2a4;
	wire			B2w2a4;
	wire			I2w2a4;
	wire			P2w2a4;
	wire			W2w2a4;
	wire			D3w2a4;
	wire			K3w2a4;
	wire			R3w2a4;
	wire			Y3w2a4;
	wire			F4w2a4;
	wire			M4w2a4;
	wire			T4w2a4;
	wire			A5w2a4;
	wire			H5w2a4;
	wire			O5w2a4;
	wire			V5w2a4;
	wire			C6w2a4;
	wire			J6w2a4;
	wire			Q6w2a4;
	wire			X6w2a4;
	wire			E7w2a4;
	wire			L7w2a4;
	wire			S7w2a4;
	wire			Z7w2a4;
	wire			G8w2a4;
	wire			N8w2a4;
	wire			U8w2a4;
	wire			B9w2a4;
	wire			I9w2a4;
	wire			P9w2a4;
	wire			W9w2a4;
	wire			Daw2a4;
	wire			Kaw2a4;
	wire			Raw2a4;
	wire			Yaw2a4;
	wire			Fbw2a4;
	wire			Mbw2a4;
	wire			Tbw2a4;
	wire			Acw2a4;
	wire			Hcw2a4;
	wire			Ocw2a4;
	wire			Vcw2a4;
	wire			Cdw2a4;
	wire			Jdw2a4;
	wire			Qdw2a4;
	wire			Xdw2a4;
	wire			Eew2a4;
	wire			Lew2a4;
	wire			Sew2a4;
	wire			Zew2a4;
	wire			Gfw2a4;
	wire			Nfw2a4;
	wire			Ufw2a4;
	wire			Bgw2a4;
	wire			Igw2a4;
	wire			Pgw2a4;
	wire			Wgw2a4;
	wire			Dhw2a4;
	wire			Khw2a4;
	wire			Rhw2a4;
	wire			Yhw2a4;
	wire			Fiw2a4;
	wire			Miw2a4;
	wire			Tiw2a4;
	wire			Ajw2a4;
	wire			Hjw2a4;
	wire			Ojw2a4;
	wire			Vjw2a4;
	wire			Ckw2a4;
	wire			Jkw2a4;
	wire			Qkw2a4;
	wire			Xkw2a4;
	wire			Elw2a4;
	wire			Llw2a4;
	wire			Slw2a4;
	wire			Zlw2a4;
	wire			Gmw2a4;
	wire			Nmw2a4;
	wire			Umw2a4;
	wire			Bnw2a4;
	wire			Inw2a4;
	wire			Pnw2a4;
	wire			Wnw2a4;
	wire			Dow2a4;
	wire			Kow2a4;
	wire			Row2a4;
	wire			Yow2a4;
	wire			Fpw2a4;
	wire			Mpw2a4;
	wire			Tpw2a4;
	wire			Aqw2a4;
	wire			Hqw2a4;
	wire			Oqw2a4;
	wire			Vqw2a4;
	wire			Crw2a4;
	wire			Jrw2a4;
	wire			Qrw2a4;
	wire			Xrw2a4;
	wire			Esw2a4;
	wire			Lsw2a4;
	wire			Ssw2a4;
	wire			Zsw2a4;
	wire			Gtw2a4;
	wire			Ntw2a4;
	wire			Utw2a4;
	wire			Buw2a4;
	wire			Iuw2a4;
	wire			Puw2a4;
	wire			Wuw2a4;
	wire			Dvw2a4;
	wire			Kvw2a4;
	wire			Rvw2a4;
	wire			Yvw2a4;
	wire			Fww2a4;
	wire			Mww2a4;
	wire			Tww2a4;
	wire			Axw2a4;
	wire			Hxw2a4;
	wire			Oxw2a4;
	wire			Vxw2a4;
	wire			Cyw2a4;
	wire			Jyw2a4;
	wire			Qyw2a4;
	wire			Xyw2a4;
	wire			Ezw2a4;
	wire			Lzw2a4;
	wire			Szw2a4;
	wire			Zzw2a4;
	wire			G0x2a4;
	wire			N0x2a4;
	wire			U0x2a4;
	wire			B1x2a4;
	wire			I1x2a4;
	wire			P1x2a4;
	wire			W1x2a4;
	wire			D2x2a4;
	wire			K2x2a4;
	wire			R2x2a4;
	wire			Y2x2a4;
	wire			F3x2a4;
	wire			M3x2a4;
	wire			T3x2a4;
	wire			A4x2a4;
	wire			H4x2a4;
	wire			O4x2a4;
	wire			V4x2a4;
	wire			C5x2a4;
	wire			J5x2a4;
	wire			Q5x2a4;
	wire			X5x2a4;
	wire			E6x2a4;
	wire			L6x2a4;
	wire			S6x2a4;
	wire			Z6x2a4;
	wire			G7x2a4;
	wire			N7x2a4;
	wire			U7x2a4;
	wire			B8x2a4;
	wire			I8x2a4;
	wire			P8x2a4;
	wire			W8x2a4;
	wire			D9x2a4;
	wire			K9x2a4;
	wire			R9x2a4;
	wire			Y9x2a4;
	wire			Fax2a4;
	wire			Max2a4;
	wire			Tax2a4;
	wire			Abx2a4;
	wire			Hbx2a4;
	wire			Obx2a4;
	wire			Vbx2a4;
	wire			Ccx2a4;
	wire			Jcx2a4;
	wire			Qcx2a4;
	wire			Xcx2a4;
	wire			Edx2a4;
	wire			Ldx2a4;
	wire			Sdx2a4;
	wire			Zdx2a4;
	wire			Gex2a4;
	wire			Nex2a4;
	wire			Uex2a4;
	wire			Bfx2a4;
	wire			Ifx2a4;
	wire			Pfx2a4;
	wire			Wfx2a4;
	wire			Dgx2a4;
	wire			Kgx2a4;
	wire			Rgx2a4;
	wire			Ygx2a4;
	wire			Fhx2a4;
	wire			Mhx2a4;
	wire			Thx2a4;
	wire			Aix2a4;
	wire			Hix2a4;
	wire			Oix2a4;
	wire			Vix2a4;
	wire			Cjx2a4;
	wire			Jjx2a4;
	wire			Qjx2a4;
	wire			Xjx2a4;
	wire			Ekx2a4;
	wire			Lkx2a4;
	wire			Skx2a4;
	wire			Zkx2a4;
	wire			Glx2a4;
	wire			Nlx2a4;
	wire			Ulx2a4;
	wire			Bmx2a4;
	wire			Imx2a4;
	wire			Pmx2a4;
	wire			Wmx2a4;
	wire			Dnx2a4;
	wire			Knx2a4;
	wire			Rnx2a4;
	wire			Ynx2a4;
	wire			Fox2a4;
	wire			Mox2a4;
	wire			Tox2a4;
	wire			Apx2a4;
	wire			Hpx2a4;
	wire			Opx2a4;
	wire			Vpx2a4;
	wire			Cqx2a4;
	wire			Jqx2a4;
	wire			Qqx2a4;
	wire			Xqx2a4;
	wire			Erx2a4;
	wire			Lrx2a4;
	wire			Srx2a4;
	wire			Zrx2a4;
	wire			Gsx2a4;
	wire			Nsx2a4;
	wire			Usx2a4;
	wire			Btx2a4;
	wire			Itx2a4;
	wire			Ptx2a4;
	wire			Wtx2a4;
	wire			Dux2a4;
	wire			Kux2a4;
	wire			Rux2a4;
	wire			Yux2a4;
	wire			Fvx2a4;
	wire			Mvx2a4;
	wire			Tvx2a4;
	wire			Awx2a4;
	wire			Hwx2a4;
	wire			Owx2a4;
	wire			Vwx2a4;
	wire			Cxx2a4;
	wire			Jxx2a4;
	wire			Qxx2a4;
	wire			Xxx2a4;
	wire			Eyx2a4;
	wire			Lyx2a4;
	wire			Syx2a4;
	wire			Zyx2a4;
	wire			Gzx2a4;
	wire			Nzx2a4;
	wire			Uzx2a4;
	wire			B0y2a4;
	wire			I0y2a4;
	wire			P0y2a4;
	wire			W0y2a4;
	wire			D1y2a4;
	wire			K1y2a4;
	wire			R1y2a4;
	wire			Y1y2a4;
	wire			F2y2a4;
	wire			M2y2a4;
	wire			T2y2a4;
	wire			A3y2a4;
	wire			H3y2a4;
	wire			O3y2a4;
	wire			V3y2a4;
	wire			C4y2a4;
	wire			J4y2a4;
	wire			Q4y2a4;
	wire			X4y2a4;
	wire			E5y2a4;
	wire			L5y2a4;
	wire			S5y2a4;
	wire			Z5y2a4;
	wire			G6y2a4;
	wire			N6y2a4;
	wire			U6y2a4;
	wire			B7y2a4;
	wire			I7y2a4;
	wire			P7y2a4;
	wire			W7y2a4;
	wire			D8y2a4;
	wire			K8y2a4;
	wire			R8y2a4;
	wire			Y8y2a4;
	wire			F9y2a4;
	wire			M9y2a4;
	wire			T9y2a4;
	wire			Aay2a4;
	wire			Hay2a4;
	wire			Oay2a4;
	wire			Vay2a4;
	wire			Cby2a4;
	wire			Jby2a4;
	wire			Qby2a4;
	wire			Xby2a4;
	wire			Ecy2a4;
	wire			Lcy2a4;
	wire			Scy2a4;
	wire			Zcy2a4;
	wire			Gdy2a4;
	wire			Ndy2a4;
	wire			Udy2a4;
	wire			Bey2a4;
	wire			Iey2a4;
	wire			Pey2a4;
	wire			Wey2a4;
	wire			Dfy2a4;
	wire			Kfy2a4;
	wire			Rfy2a4;
	wire			Yfy2a4;
	wire			Fgy2a4;
	wire			Mgy2a4;
	wire			Tgy2a4;
	wire			Ahy2a4;
	wire			Hhy2a4;
	wire			Ohy2a4;
	wire			Vhy2a4;
	wire			Ciy2a4;
	wire			Jiy2a4;
	wire			Qiy2a4;
	wire			Xiy2a4;
	wire			Ejy2a4;
	wire			Ljy2a4;
	wire			Sjy2a4;
	wire			Zjy2a4;
	wire			Gky2a4;
	wire			Nky2a4;
	wire			Uky2a4;
	wire			Bly2a4;
	wire			Ily2a4;
	wire			Ply2a4;
	wire			Wly2a4;
	wire			Dmy2a4;
	wire			Kmy2a4;
	wire			Rmy2a4;
	wire			Ymy2a4;
	wire			Fny2a4;
	wire			Mny2a4;
	wire			Tny2a4;
	wire			Aoy2a4;
	wire			Hoy2a4;
	wire			Ooy2a4;
	wire			Voy2a4;
	wire			Cpy2a4;
	wire			Jpy2a4;
	wire			Qpy2a4;
	wire			Xpy2a4;
	wire			Eqy2a4;
	wire			Lqy2a4;
	wire			Sqy2a4;
	wire			Zqy2a4;
	wire			Gry2a4;
	wire			Nry2a4;
	wire			Ury2a4;
	wire			Bsy2a4;
	wire			Isy2a4;
	wire			Psy2a4;
	wire			Wsy2a4;
	wire			Dty2a4;
	wire			Kty2a4;
	wire			Rty2a4;
	wire			Yty2a4;
	wire			Fuy2a4;
	wire			Muy2a4;
	wire			Tuy2a4;
	wire			Avy2a4;
	wire			Hvy2a4;
	wire			Ovy2a4;
	wire			Vvy2a4;
	wire			Cwy2a4;
	wire			Jwy2a4;
	wire			Qwy2a4;
	wire			Xwy2a4;
	wire			Exy2a4;
	wire			Lxy2a4;
	wire			Sxy2a4;
	wire			Zxy2a4;
	wire			Gyy2a4;
	wire			Nyy2a4;
	wire			Uyy2a4;
	wire			Bzy2a4;
	wire			Izy2a4;
	wire			Pzy2a4;
	wire			Wzy2a4;
	wire			D0z2a4;
	wire			K0z2a4;
	wire			R0z2a4;
	wire			Y0z2a4;
	wire			F1z2a4;
	wire			M1z2a4;
	wire			T1z2a4;
	wire			A2z2a4;
	wire			H2z2a4;
	wire			O2z2a4;
	wire			V2z2a4;
	wire			C3z2a4;
	wire			J3z2a4;
	wire			Q3z2a4;
	wire			X3z2a4;
	wire			E4z2a4;
	wire			L4z2a4;
	wire			S4z2a4;
	wire			Z4z2a4;
	wire			G5z2a4;
	wire			N5z2a4;
	wire			U5z2a4;
	wire			B6z2a4;
	wire			I6z2a4;
	wire			P6z2a4;
	wire			W6z2a4;
	wire			D7z2a4;
	wire			K7z2a4;
	wire			R7z2a4;
	wire			Y7z2a4;
	wire			F8z2a4;
	wire			M8z2a4;
	wire			T8z2a4;
	wire			A9z2a4;
	wire			H9z2a4;
	wire			O9z2a4;
	wire			V9z2a4;
	wire			Caz2a4;
	wire			Jaz2a4;
	wire			Qaz2a4;
	wire			Xaz2a4;
	wire			Ebz2a4;
	wire			Lbz2a4;
	wire			Sbz2a4;
	wire			Zbz2a4;
	wire			Gcz2a4;
	wire			Ncz2a4;
	wire			Ucz2a4;
	wire			Bdz2a4;
	wire			Idz2a4;
	wire			Pdz2a4;
	wire			Wdz2a4;
	wire			Dez2a4;
	wire			Kez2a4;
	wire			Rez2a4;
	wire			Yez2a4;
	wire			Ffz2a4;
	wire			Mfz2a4;
	wire			Tfz2a4;
	wire			Agz2a4;
	wire			Hgz2a4;
	wire			Ogz2a4;
	wire			Vgz2a4;
	wire			Chz2a4;
	wire			Jhz2a4;
	wire			Qhz2a4;
	wire			Xhz2a4;
	wire			Eiz2a4;
	wire			Liz2a4;
	wire			Siz2a4;
	wire			Ziz2a4;
	wire			Gjz2a4;
	wire			Njz2a4;
	wire			Ujz2a4;
	wire			Bkz2a4;
	wire			Ikz2a4;
	wire			Pkz2a4;
	wire			Wkz2a4;
	wire			Dlz2a4;
	wire			Klz2a4;
	wire			Rlz2a4;
	wire			Ylz2a4;
	wire			Fmz2a4;
	wire			Mmz2a4;
	wire			Tmz2a4;
	wire			Anz2a4;
	wire			Hnz2a4;
	wire			Onz2a4;
	wire			Vnz2a4;
	wire			Coz2a4;
	wire			Joz2a4;
	wire			Qoz2a4;
	wire			Xoz2a4;
	wire			Epz2a4;
	wire			Lpz2a4;
	wire			Spz2a4;
	wire			Zpz2a4;
	wire			Gqz2a4;
	wire			Nqz2a4;
	wire			Uqz2a4;
	wire			Brz2a4;
	wire			Irz2a4;
	wire			Prz2a4;
	wire			Wrz2a4;
	wire			Dsz2a4;
	wire			Ksz2a4;
	wire			Rsz2a4;
	wire			Ysz2a4;
	wire			Ftz2a4;
	wire			Mtz2a4;
	wire			Ttz2a4;
	wire			Auz2a4;
	wire			Huz2a4;
	wire			Ouz2a4;
	wire			Vuz2a4;
	wire			Cvz2a4;
	wire			Jvz2a4;
	wire			Qvz2a4;
	wire			Xvz2a4;
	wire			Ewz2a4;
	wire			Lwz2a4;
	wire			Swz2a4;
	wire			Zwz2a4;
	wire			Gxz2a4;
	wire			Nxz2a4;
	wire			Uxz2a4;
	wire			Byz2a4;
	wire			Iyz2a4;
	wire			Pyz2a4;
	wire			Wyz2a4;
	wire			Dzz2a4;
	wire			Kzz2a4;
	wire			Rzz2a4;
	wire			Yzz2a4;
	wire			F003a4;
	wire			M003a4;
	wire			T003a4;
	wire			A103a4;
	wire			H103a4;
	wire			O103a4;
	wire			V103a4;
	wire			C203a4;
	wire			J203a4;
	wire			Q203a4;
	wire			X203a4;
	wire			E303a4;
	wire			L303a4;
	wire			S303a4;
	wire			Z303a4;
	wire			G403a4;
	wire			N403a4;
	wire			U403a4;
	wire			B503a4;
	wire			I503a4;
	wire			P503a4;
	wire			W503a4;
	wire			D603a4;
	wire			K603a4;
	wire			R603a4;
	wire			Y603a4;
	wire			F703a4;
	wire			M703a4;
	wire			T703a4;
	wire			A803a4;
	wire			H803a4;
	wire			O803a4;
	wire			V803a4;
	wire			C903a4;
	wire			J903a4;
	wire			Q903a4;
	wire			X903a4;
	wire			Ea03a4;
	wire			La03a4;
	wire			Sa03a4;
	wire			Za03a4;
	wire			Gb03a4;
	wire			Nb03a4;
	wire			Ub03a4;
	wire			Bc03a4;
	wire			Ic03a4;
	wire			Pc03a4;
	wire			Wc03a4;
	wire			Dd03a4;
	wire			Kd03a4;
	wire			Rd03a4;
	wire			Yd03a4;
	wire			Fe03a4;
	wire			Me03a4;
	wire			Te03a4;
	wire			Af03a4;
	wire			Hf03a4;
	wire			Of03a4;
	wire			Vf03a4;
	wire			Cg03a4;
	wire			Jg03a4;
	wire			Qg03a4;
	wire			Xg03a4;
	wire			Eh03a4;
	wire			Lh03a4;
	wire			Sh03a4;
	wire			Zh03a4;
	wire			Gi03a4;
	wire			Ni03a4;
	wire			Ui03a4;
	wire			Bj03a4;
	wire			Ij03a4;
	wire			Pj03a4;
	wire			Wj03a4;
	wire			Dk03a4;
	wire			Kk03a4;
	wire			Rk03a4;
	wire			Yk03a4;
	wire			Fl03a4;
	wire			Ml03a4;
	wire			Tl03a4;
	wire			Am03a4;
	wire			Hm03a4;
	wire			Om03a4;
	wire			Vm03a4;
	wire			Cn03a4;
	wire			Jn03a4;
	wire			Qn03a4;
	wire			Xn03a4;
	wire			Eo03a4;
	wire			Lo03a4;
	wire			So03a4;
	wire			Zo03a4;
	wire			Gp03a4;
	wire			Np03a4;
	wire			Up03a4;
	wire			Bq03a4;
	wire			Iq03a4;
	wire			Pq03a4;
	wire			Wq03a4;
	wire			Dr03a4;
	wire			Kr03a4;
	wire			Rr03a4;
	wire			Yr03a4;
	wire			Fs03a4;
	wire			Ms03a4;
	wire			Ts03a4;
	wire			At03a4;
	wire			Ht03a4;
	wire			Ot03a4;
	wire			Vt03a4;
	wire			Cu03a4;
	wire			Ju03a4;
	wire			Qu03a4;
	wire			Xu03a4;
	wire			Ev03a4;
	wire			Lv03a4;
	wire			Sv03a4;
	wire			Zv03a4;
	wire			Gw03a4;
	wire			Nw03a4;
	wire			Uw03a4;
	wire			Bx03a4;
	wire			Ix03a4;
	wire			Px03a4;
	wire			Wx03a4;
	wire			Dy03a4;
	wire			Ky03a4;
	wire			Ry03a4;
	wire			Yy03a4;
	wire			Fz03a4;
	wire			Mz03a4;
	wire			Tz03a4;
	wire			A013a4;
	wire			H013a4;
	wire			O013a4;
	wire			V013a4;
	wire			C113a4;
	wire			J113a4;
	wire			Q113a4;
	wire			X113a4;
	wire			E213a4;
	wire			L213a4;
	wire			S213a4;
	wire			Z213a4;
	wire			G313a4;
	wire			N313a4;
	wire			U313a4;
	wire			B413a4;
	wire			I413a4;
	wire			P413a4;
	wire			W413a4;
	wire			D513a4;
	wire			K513a4;
	wire			R513a4;
	wire			Y513a4;
	wire			F613a4;
	wire			M613a4;
	wire			T613a4;
	wire			A713a4;
	wire			H713a4;
	wire			O713a4;
	wire			V713a4;
	wire			C813a4;
	wire			J813a4;
	wire			Q813a4;
	wire			X813a4;
	wire			E913a4;
	wire			L913a4;
	wire			S913a4;
	wire			Z913a4;
	wire			Ga13a4;
	wire			Na13a4;
	wire			Ua13a4;
	wire			Bb13a4;
	wire			Ib13a4;
	wire			Pb13a4;
	wire			Wb13a4;
	wire			Dc13a4;
	wire			Kc13a4;
	wire			Rc13a4;
	wire			Yc13a4;
	wire			Fd13a4;
	wire			Md13a4;
	wire			Td13a4;
	wire			Ae13a4;
	wire			He13a4;
	wire			Oe13a4;
	wire			Ve13a4;
	wire			Cf13a4;
	wire			Jf13a4;
	wire			Qf13a4;
	wire			Xf13a4;
	wire			Eg13a4;
	wire			Lg13a4;
	wire			Sg13a4;
	wire			Zg13a4;
	wire			Gh13a4;
	wire			Nh13a4;
	wire			Uh13a4;
	wire			Bi13a4;
	wire			Ii13a4;
	wire			Pi13a4;
	wire			Wi13a4;
	wire			Dj13a4;
	wire			Kj13a4;
	wire			Rj13a4;
	wire			Yj13a4;
	wire			Fk13a4;
	wire			Mk13a4;
	wire			Tk13a4;
	wire			Al13a4;
	wire			Hl13a4;
	wire			Ol13a4;
	wire			Vl13a4;
	wire			Cm13a4;
	wire			Jm13a4;
	wire			Qm13a4;
	wire			Xm13a4;
	wire			En13a4;
	wire			Ln13a4;
	wire			Sn13a4;
	wire			Zn13a4;
	wire			Go13a4;
	wire			No13a4;
	wire			Uo13a4;
	wire			Bp13a4;
	wire			Ip13a4;
	wire			Pp13a4;
	wire			Wp13a4;
	wire			Dq13a4;
	wire			Kq13a4;
	wire			Rq13a4;
	wire			Yq13a4;
	wire			Fr13a4;
	wire			Mr13a4;
	wire			Tr13a4;
	wire			As13a4;
	wire			Hs13a4;
	wire			Os13a4;
	wire			Vs13a4;
	wire			Ct13a4;
	wire			Jt13a4;
	wire			Qt13a4;
	wire			Xt13a4;
	wire			Eu13a4;
	wire			Lu13a4;
	wire			Su13a4;
	wire			Zu13a4;
	wire			Gv13a4;
	wire			Nv13a4;
	wire			Uv13a4;
	wire			Bw13a4;
	wire			Iw13a4;
	wire			Pw13a4;
	wire			Ww13a4;
	wire			Dx13a4;
	wire			Kx13a4;
	wire			Rx13a4;
	wire			Yx13a4;
	wire			Fy13a4;
	wire			My13a4;
	wire			Ty13a4;
	wire			Az13a4;
	wire			Hz13a4;
	wire			Oz13a4;
	wire			Vz13a4;
	wire			C023a4;
	wire			J023a4;
	wire			Q023a4;
	wire			X023a4;
	wire			E123a4;
	wire			L123a4;
	wire			S123a4;
	wire			Z123a4;
	wire			G223a4;
	wire			N223a4;
	wire			U223a4;
	wire			B323a4;
	wire			I323a4;
	wire			P323a4;
	wire			W323a4;
	wire			D423a4;
	wire			K423a4;
	wire			R423a4;
	wire			Y423a4;
	wire			F523a4;
	wire			M523a4;
	wire			T523a4;
	wire			A623a4;
	wire			H623a4;
	wire			O623a4;
	wire			V623a4;
	wire			C723a4;
	wire			J723a4;
	wire			Q723a4;
	wire			X723a4;
	wire			E823a4;
	wire			L823a4;
	wire			S823a4;
	wire			Z823a4;
	wire			G923a4;
	wire			N923a4;
	wire			U923a4;
	wire			Ba23a4;
	wire			Ia23a4;
	wire			Pa23a4;
	wire			Wa23a4;
	wire			Db23a4;
	wire			Kb23a4;
	wire			Rb23a4;
	wire			Yb23a4;
	wire			Fc23a4;
	wire			Mc23a4;
	wire			Tc23a4;
	wire			Ad23a4;
	wire			Hd23a4;
	wire			Od23a4;
	wire			Vd23a4;
	wire			Ce23a4;
	wire			Je23a4;
	wire			Qe23a4;
	wire			Xe23a4;
	wire			Ef23a4;
	wire			Lf23a4;
	wire			Sf23a4;
	wire			Zf23a4;
	wire			Gg23a4;
	wire			Ng23a4;
	wire			Ug23a4;
	wire			Bh23a4;
	wire			Ih23a4;
	wire			Ph23a4;
	wire			Wh23a4;
	wire			Di23a4;
	wire			Ki23a4;
	wire			Ri23a4;
	wire			Yi23a4;
	wire			Fj23a4;
	wire			Mj23a4;
	wire			Tj23a4;
	wire			Ak23a4;
	wire			Hk23a4;
	wire			Ok23a4;
	wire			Vk23a4;
	wire			Cl23a4;
	wire			Jl23a4;
	wire			Ql23a4;
	wire			Xl23a4;
	wire			Em23a4;
	wire			Lm23a4;
	wire			Sm23a4;
	wire			Zm23a4;
	wire			Gn23a4;
	wire			Nn23a4;
	wire			Un23a4;
	wire			Bo23a4;
	wire			Io23a4;
	wire			Po23a4;
	wire			Wo23a4;
	wire			Dp23a4;
	wire			Kp23a4;
	wire			Rp23a4;
	wire			Yp23a4;
	wire			Fq23a4;
	wire			Mq23a4;
	wire			Tq23a4;
	wire			Ar23a4;
	wire			Hr23a4;
	wire			Or23a4;
	wire			Vr23a4;
	wire			Cs23a4;
	wire			Js23a4;
	wire			Qs23a4;
	wire			Xs23a4;
	wire			Et23a4;
	wire			Lt23a4;
	wire			St23a4;
	wire			Zt23a4;
	wire			Gu23a4;
	wire			Nu23a4;
	wire			Uu23a4;
	wire			Bv23a4;
	wire			Iv23a4;
	wire			Pv23a4;
	wire			Wv23a4;
	wire			Dw23a4;
	wire			Kw23a4;
	wire			Rw23a4;
	wire			Yw23a4;
	wire			Fx23a4;
	wire			Mx23a4;
	wire			Tx23a4;
	wire			Ay23a4;
	wire			Hy23a4;
	wire			Oy23a4;
	wire			Vy23a4;
	wire			Cz23a4;
	wire			Jz23a4;
	wire			Qz23a4;
	wire			Xz23a4;
	wire			E033a4;
	wire			L033a4;
	wire			S033a4;
	wire			Z033a4;
	wire			G133a4;
	wire			N133a4;
	wire			U133a4;
	wire			B233a4;
	wire			I233a4;
	wire			P233a4;
	wire			W233a4;
	wire			D333a4;
	wire			K333a4;
	wire			R333a4;
	wire			Y333a4;
	wire			F433a4;
	wire			M433a4;
	wire			T433a4;
	wire			A533a4;
	wire			H533a4;
	wire			O533a4;
	wire			V533a4;
	wire			C633a4;
	wire			J633a4;
	wire			Q633a4;
	wire			X633a4;
	wire			E733a4;
	wire			L733a4;
	wire			S733a4;
	wire			Z733a4;
	wire			G833a4;
	wire			N833a4;
	wire			U833a4;
	wire			B933a4;
	wire			I933a4;
	wire			P933a4;
	wire			W933a4;
	wire			Da33a4;
	wire			Ka33a4;
	wire			Ra33a4;
	wire			Ya33a4;
	wire			Fb33a4;
	wire			Mb33a4;
	wire			Tb33a4;
	wire			Ac33a4;
	wire			Hc33a4;
	wire			Oc33a4;
	wire			Vc33a4;
	wire			Cd33a4;
	wire			Jd33a4;
	wire			Qd33a4;
	wire			Xd33a4;
	wire			Ee33a4;
	wire			Le33a4;
	wire			Se33a4;
	wire			Ze33a4;
	wire			Gf33a4;
	wire			Nf33a4;
	wire			Uf33a4;
	wire			Bg33a4;
	wire			Ig33a4;
	wire			Pg33a4;
	wire			Wg33a4;
	wire			Dh33a4;
	wire			Kh33a4;
	wire			Rh33a4;
	wire			Yh33a4;
	wire			Fi33a4;
	wire			Mi33a4;
	wire			Ti33a4;
	wire			Aj33a4;
	wire			Hj33a4;
	wire			Oj33a4;
	wire			Vj33a4;
	wire			Ck33a4;
	wire			Jk33a4;
	wire			Qk33a4;
	wire			Xk33a4;
	wire			El33a4;
	wire			Ll33a4;
	wire			Sl33a4;
	wire			Zl33a4;
	wire			Gm33a4;
	wire			Nm33a4;
	wire			Um33a4;
	wire			Bn33a4;
	wire			In33a4;
	wire			Pn33a4;
	wire			Wn33a4;
	wire			Do33a4;
	wire			Ko33a4;
	wire			Ro33a4;
	wire			Yo33a4;
	wire			Fp33a4;
	wire			Mp33a4;
	wire			Tp33a4;
	wire			Aq33a4;
	wire			Hq33a4;
	wire			Oq33a4;
	wire			Vq33a4;
	wire			Cr33a4;
	wire			Jr33a4;
	wire			Qr33a4;
	wire			Xr33a4;
	wire			Es33a4;
	wire			Ls33a4;
	wire			Ss33a4;
	wire			Zs33a4;
	wire			Gt33a4;
	wire			Nt33a4;
	wire			Ut33a4;
	wire			Bu33a4;
	wire			Iu33a4;
	wire			Pu33a4;
	wire			Wu33a4;
	wire			Dv33a4;
	wire			Kv33a4;
	wire			Rv33a4;
	wire			Yv33a4;
	wire			Fw33a4;
	wire			Mw33a4;
	wire			Tw33a4;
	wire			Ax33a4;
	wire			Hx33a4;
	wire			Ox33a4;
	wire			Vx33a4;
	wire			Cy33a4;
	wire			Jy33a4;
	wire			Qy33a4;
	wire			Xy33a4;
	wire			Ez33a4;
	wire			Lz33a4;
	wire			Sz33a4;
	wire			Zz33a4;
	wire			G043a4;
	wire			N043a4;
	wire			U043a4;
	wire			B143a4;
	wire			I143a4;
	wire			P143a4;
	wire			W143a4;
	wire			D243a4;
	wire			K243a4;
	wire			R243a4;
	wire			Y243a4;
	wire			F343a4;
	wire			M343a4;
	wire			T343a4;
	wire			A443a4;
	wire			H443a4;
	wire			O443a4;
	wire			V443a4;
	wire			C543a4;
	wire			J543a4;
	wire			Q543a4;
	wire			X543a4;
	wire			E643a4;
	wire			L643a4;
	wire			S643a4;
	wire			Z643a4;
	wire			G743a4;
	wire			N743a4;
	wire			U743a4;
	wire			B843a4;
	wire			I843a4;
	wire			P843a4;
	wire			W843a4;
	wire			D943a4;
	wire			K943a4;
	wire			R943a4;
	wire			Y943a4;
	wire			Fa43a4;
	wire			Ma43a4;
	wire			Ta43a4;
	wire			Ab43a4;
	wire			Hb43a4;
	wire			Ob43a4;
	wire			Vb43a4;
	wire			Cc43a4;
	wire			Jc43a4;
	wire			Qc43a4;
	wire			Xc43a4;
	wire			Ed43a4;
	wire			Ld43a4;
	wire			Sd43a4;
	wire			Zd43a4;
	wire			Ge43a4;
	wire			Ne43a4;
	wire			Ue43a4;
	wire			Bf43a4;
	wire			If43a4;
	wire			Pf43a4;
	wire			Wf43a4;
	wire			Dg43a4;
	wire			Kg43a4;
	wire			Rg43a4;
	wire			Yg43a4;
	wire			Fh43a4;
	wire			Mh43a4;
	wire			Th43a4;
	wire			Ai43a4;
	wire			Hi43a4;
	wire			Oi43a4;
	wire			Vi43a4;
	wire			Cj43a4;
	wire			Jj43a4;
	wire			Qj43a4;
	wire			Xj43a4;
	wire			Ek43a4;
	wire			Lk43a4;
	wire			Sk43a4;
	wire			Zk43a4;
	wire			Gl43a4;
	wire			Nl43a4;
	wire			Ul43a4;
	wire			Bm43a4;
	wire			Im43a4;
	wire			Pm43a4;
	wire			Wm43a4;
	wire			Dn43a4;
	wire			Kn43a4;
	wire			Rn43a4;
	wire			Yn43a4;
	wire			Fo43a4;
	wire			Mo43a4;
	wire			To43a4;
	wire			Ap43a4;
	wire			Hp43a4;
	wire			Op43a4;
	wire			Vp43a4;
	wire			Cq43a4;
	wire			Jq43a4;
	wire			Qq43a4;
	wire			Xq43a4;
	wire			Er43a4;
	wire			Lr43a4;
	wire			Sr43a4;
	wire			Zr43a4;
	wire			Gs43a4;
	wire			Ns43a4;
	wire			Us43a4;
	wire			Bt43a4;
	wire			It43a4;
	wire			Pt43a4;
	wire			Wt43a4;
	wire			Du43a4;
	wire			Ku43a4;
	wire			Ru43a4;
	wire			Yu43a4;
	wire			Fv43a4;
	wire			Mv43a4;
	wire			Tv43a4;
	wire			Aw43a4;
	wire			Hw43a4;
	wire			Ow43a4;
	wire			Vw43a4;
	wire			Cx43a4;
	wire			Jx43a4;
	wire			Qx43a4;
	wire			Xx43a4;
	wire			Ey43a4;
	wire			Ly43a4;
	wire			Sy43a4;
	wire			Zy43a4;
	wire			Gz43a4;
	wire			Nz43a4;
	wire			Uz43a4;
	wire			B053a4;
	wire			I053a4;
	wire			P053a4;
	wire			W053a4;
	wire			D153a4;
	wire			K153a4;
	wire			R153a4;
	wire			Y153a4;
	wire			F253a4;
	wire			M253a4;
	wire			T253a4;
	wire			A353a4;
	wire			H353a4;
	wire			O353a4;
	wire			V353a4;
	wire			C453a4;
	wire			J453a4;
	wire			Q453a4;
	wire			X453a4;
	wire			E553a4;
	wire			L553a4;
	wire			S553a4;
	wire			Z553a4;
	wire			G653a4;
	wire			N653a4;
	wire			U653a4;
	wire			B753a4;
	wire			I753a4;
	wire			P753a4;
	wire			W753a4;
	wire			D853a4;
	wire			K853a4;
	wire			R853a4;
	wire			Y853a4;
	wire			F953a4;
	wire			M953a4;
	wire			T953a4;
	wire			Aa53a4;
	wire			Ha53a4;
	wire			Oa53a4;
	wire			Va53a4;
	wire			Cb53a4;
	wire			Jb53a4;
	wire			Qb53a4;
	wire			Xb53a4;
	wire			Ec53a4;
	wire			Lc53a4;
	wire			Sc53a4;
	wire			Zc53a4;
	wire			Gd53a4;
	wire			Nd53a4;
	wire			Ud53a4;
	wire			Be53a4;
	wire			Ie53a4;
	wire			Pe53a4;
	wire			We53a4;
	wire			Df53a4;
	wire			Kf53a4;
	wire			Rf53a4;
	wire			Yf53a4;
	wire			Fg53a4;
	wire			Mg53a4;
	wire			Tg53a4;
	wire			Ah53a4;
	wire			Hh53a4;
	wire			Oh53a4;
	wire			Vh53a4;
	wire			Ci53a4;
	wire			Ji53a4;
	wire			Qi53a4;
	wire			Xi53a4;
	wire			Ej53a4;
	wire			Lj53a4;
	wire			Sj53a4;
	wire			Zj53a4;
	wire			Gk53a4;
	wire			Nk53a4;
	wire			Uk53a4;
	wire			Bl53a4;
	wire			Il53a4;
	wire			Pl53a4;
	wire			Wl53a4;
	wire			Dm53a4;
	wire			Km53a4;
	wire			Rm53a4;
	wire			Ym53a4;
	wire			Fn53a4;
	wire			Mn53a4;
	wire			Tn53a4;
	wire			Ao53a4;
	wire			Ho53a4;
	wire			Oo53a4;
	wire			Vo53a4;
	wire			Cp53a4;
	wire			Jp53a4;
	wire			Qp53a4;
	wire			Xp53a4;
	wire			Eq53a4;
	wire			Lq53a4;
	wire			Sq53a4;
	wire			Zq53a4;
	wire			Gr53a4;
	wire			Nr53a4;
	wire			Ur53a4;
	wire			Bs53a4;
	wire			Is53a4;
	wire			Ps53a4;
	wire			Ws53a4;
	wire			Dt53a4;
	wire			Kt53a4;
	wire			Rt53a4;
	wire			Yt53a4;
	wire			Fu53a4;
	wire			Mu53a4;
	wire			Tu53a4;
	wire			Av53a4;
	wire			Hv53a4;
	wire			Ov53a4;
	wire			Vv53a4;
	wire			Cw53a4;
	wire			Jw53a4;
	wire			Qw53a4;
	wire			Xw53a4;
	wire			Ex53a4;
	wire			Lx53a4;
	wire			Sx53a4;
	wire			Zx53a4;
	wire			Gy53a4;
	wire			Ny53a4;
	wire			Uy53a4;
	wire			Bz53a4;
	wire			Iz53a4;
	wire			Pz53a4;
	wire			Wz53a4;
	wire			D063a4;
	wire			K063a4;
	wire			R063a4;
	wire			Y063a4;
	wire			F163a4;
	wire			M163a4;
	wire			T163a4;
	wire			A263a4;
	wire			H263a4;
	wire			O263a4;
	wire			V263a4;
	wire			C363a4;
	wire			J363a4;
	wire			Q363a4;
	wire			X363a4;
	wire			E463a4;
	wire			L463a4;
	wire			S463a4;
	wire			Z463a4;
	wire			G563a4;
	wire			N563a4;
	wire			U563a4;
	wire			B663a4;
	wire			I663a4;
	wire			P663a4;
	wire			W663a4;
	wire			D763a4;
	wire			K763a4;
	wire			R763a4;
	wire			Y763a4;
	wire			F863a4;
	wire			M863a4;
	wire			T863a4;
	wire			A963a4;
	wire			H963a4;
	wire			O963a4;
	wire			V963a4;
	wire			Ca63a4;
	wire			Ja63a4;
	wire			Qa63a4;
	wire			Xa63a4;
	wire			Eb63a4;
	wire			Lb63a4;
	wire			Sb63a4;
	wire			Zb63a4;
	wire			Gc63a4;
	wire			Nc63a4;
	wire			Uc63a4;
	wire			Bd63a4;
	wire			Id63a4;
	wire			Pd63a4;
	wire			Wd63a4;
	wire			De63a4;
	wire			Ke63a4;
	wire			Re63a4;
	wire			Ye63a4;
	wire			Ff63a4;
	wire			Mf63a4;
	wire			Tf63a4;
	wire			Ag63a4;
	wire			Hg63a4;
	wire			Og63a4;
	wire			Vg63a4;
	wire			Ch63a4;
	wire			Jh63a4;
	wire			Qh63a4;
	wire			Xh63a4;
	wire			Ei63a4;
	wire			Li63a4;
	wire			Si63a4;
	wire			Zi63a4;
	wire			Gj63a4;
	wire	[5:0]		Nj63a4;
	wire	[30:0]		Tk63a4;
	wire	[3:0]		Km63a4;
	wire	[30:2]		Ao63a4;
	wire	[31:0]		Qp63a4;
	wire	[30:0]		Cr63a4;
	wire	[1:0]		Vs63a4;
	wire	[23:0]		Pu63a4;
	wire	[1:0]		Hw63a4;
	wire	[1:0]		Xx63a4;
	wire	[7:0]		Nz63a4;
	wire	[23:0]		H173a4;
	wire	[1:0]		D373a4;
	wire	[23:0]		X473a4;
	wire	[3:0]		R673a4;
	wire	[3:0]		K873a4;
	wire			Fa73a4;
	reg			Db73a4;
	reg			Ed73a4;
	reg			Cf73a4;
	reg			Bh73a4;
	reg			Aj73a4;
	reg			Yk73a4;
	reg			Um73a4;
	reg			Xo73a4;
	reg			Wq73a4;
	reg			Ws73a4;
	reg			Qu73a4;
	reg			Lw73a4;
	reg			Fy73a4;
	reg			F083a4;
	reg			F283a4;
	reg			F483a4;
	reg			B683a4;
	reg			A883a4;
	reg			Z983a4;
	reg			Yb83a4;
	reg			Vd83a4;
	reg			Vf83a4;
	reg			Vh83a4;
	reg			Vj83a4;
	reg			Vl83a4;
	reg			Vn83a4;
	reg			Sp83a4;
	reg			Rr83a4;
	reg			Nt83a4;
	reg			Kv83a4;
	reg			Hx83a4;
	reg			Gz83a4;
	reg			F193a4;
	reg			I393a4;
	reg			H593a4;
	reg			G793a4;
	reg			E993a4;
	reg			Cb93a4;
	reg			Ad93a4;
	reg			Ve93a4;
	reg			Rg93a4;
	reg			Qi93a4;
	reg			Pk93a4;
	reg			Om93a4;
	reg			Lo93a4;
	reg			Lq93a4;
	reg			Ms93a4;
	reg			Mu93a4;
	reg			Nw93a4;
	reg			Ly93a4;
	reg			J0a3a4;
	reg			H2a3a4;
	reg			D4a3a4;
	reg			Z5a3a4;
	reg			B8a3a4;
	reg			Daa3a4;
	reg			Cca3a4;
	reg			Bea3a4;
	reg			Yfa3a4;
	reg			Yha3a4;
	reg			Aka3a4;
	reg			Cma3a4;
	reg			Boa3a4;
	reg			Upa3a4;
	reg			Tra3a4;
	reg			Pta3a4;
	reg			Mva3a4;
	reg			Mxa3a4;
	reg			Oza3a4;
	reg			Q1b3a4;
	reg			N3b3a4;
	reg			N5b3a4;
	reg			P7b3a4;
	reg			R9b3a4;
	reg			Rbb3a4;
	reg			Rdb3a4;
	reg			Lfb3a4;
	reg			Lhb3a4;
	reg			Ljb3a4;
	reg			Ilb3a4;
	reg			Dnb3a4;
	reg			Cpb3a4;
	reg			Crb3a4;
	reg			Ctb3a4;
	reg			Dvb3a4;
	reg			Axb3a4;
	reg			Azb3a4;
	reg			A1c3a4;
	reg			A3c3a4;
	reg			X4c3a4;
	reg			X6c3a4;
	reg			Z8c3a4;
	reg			Bbc3a4;
	reg			Ddc3a4;
	reg			Cfc3a4;
	reg			Bhc3a4;
	reg			Cjc3a4;
	reg			Blc3a4;
	reg			Anc3a4;
	reg			Yoc3a4;
	reg			Brc3a4;
	reg			Atc3a4;
	reg			Xuc3a4;
	reg			Xwc3a4;
	reg			Zyc3a4;
	reg			B1d3a4;
	reg			X2d3a4;
	reg			X4d3a4;
	reg			X6d3a4;
	reg			X8d3a4;
	reg			Yad3a4;
	reg			Xcd3a4;
	reg			Zed3a4;
	reg			Bhd3a4;
	reg			Yid3a4;
	reg			Ykd3a4;
	reg			Ymd3a4;
	reg			Yod3a4;
	reg			Vqd3a4;
	reg			Vsd3a4;
	reg			Wud3a4;
	reg			Swd3a4;
	reg			Ryd3a4;
	reg			S0e3a4;
	reg			P2e3a4;
	reg			P4e3a4;
	reg			P6e3a4;
	reg			P8e3a4;
	reg			Mae3a4;
	reg			Mce3a4;
	reg			Lee3a4;
	reg			Kge3a4;
	reg			Iie3a4;
	reg			Hke3a4;
	reg			Fme3a4;
	reg			Doe3a4;
	reg			Zpe3a4;
	reg			Vre3a4;
	reg			Rte3a4;
	reg			Pve3a4;
	reg			Jxe3a4;
	reg			Jze3a4;
	reg			G1f3a4;
	reg			G3f3a4;
	reg			G5f3a4;
	reg			F7f3a4;
	reg			E9f3a4;
	reg			Dbf3a4;
	reg			Adf3a4;
	reg			Xef3a4;
	reg			Xgf3a4;
	reg			Xif3a4;
	reg			Xkf3a4;
	reg			Umf3a4;
	reg			Uof3a4;
	reg			Uqf3a4;
	reg			Usf3a4;
	reg			Quf3a4;
	reg			Rwf3a4;
	reg			Oyf3a4;
	reg			N0g3a4;
	reg			M2g3a4;
	reg			L4g3a4;
	reg			I6g3a4;
	reg			I8g3a4;
	reg			Iag3a4;
	reg			Icg3a4;
	reg			Heg3a4;
	reg			Hgg3a4;
	reg			Jig3a4;
	reg			Ikg3a4;
	reg			Hmg3a4;
	reg			Gog3a4;
	reg			Dqg3a4;
	reg			Csg3a4;
	reg			Cug3a4;
	reg			Cwg3a4;
	reg			Cyg3a4;
	reg			C0h3a4;
	reg			C2h3a4;
	reg			C4h3a4;
	reg			B6h3a4;
	reg			A8h3a4;
	reg			Z9h3a4;
	reg			Ybh3a4;
	reg			Xdh3a4;
	reg			Wfh3a4;
	reg			Vhh3a4;
	reg			Ujh3a4;
	reg			Tlh3a4;
	reg			Snh3a4;
	reg			Sph3a4;
	reg			Orh3a4;
	reg			Kth3a4;
	reg			Gvh3a4;
	reg			Cxh3a4;
	reg			Yyh3a4;
	reg			V0i3a4;
	reg			R2i3a4;
	reg			O4i3a4;
	reg			L6i3a4;
	reg			I8i3a4;
	reg			Iai3a4;
	reg			Hci3a4;
	reg			Gei3a4;
	reg			Fgi3a4;
	reg			Eii3a4;
	reg			Eki3a4;
	reg			Emi3a4;
	reg			Eoi3a4;
	reg			Eqi3a4;
	reg			Esi3a4;
	reg			Eui3a4;
	reg			Dwi3a4;
	reg			Cyi3a4;
	reg			Zzi3a4;
	reg			Y1j3a4;
	reg			X3j3a4;
	reg			W5j3a4;
	reg			V7j3a4;
	reg			U9j3a4;
	reg			Ubj3a4;
	reg			Udj3a4;
	reg			Ufj3a4;
	reg			Rhj3a4;
	reg			Rjj3a4;
	reg			Qlj3a4;
	reg			Qnj3a4;
	reg			Tpj3a4;
	reg			Srj3a4;
	reg			Rtj3a4;
	reg			Qvj3a4;
	reg			Pxj3a4;
	reg			Ozj3a4;
	reg			N1k3a4;
	reg			M3k3a4;
	reg			M5k3a4;
	reg			L7k3a4;
	reg			K9k3a4;
	reg			Jbk3a4;
	reg			Idk3a4;
	reg			Hfk3a4;
	reg			Ghk3a4;
	reg			Fjk3a4;
	reg			Flk3a4;
	reg			Fnk3a4;
	reg			Fpk3a4;
	reg			Frk3a4;
	reg			Ftk3a4;
	reg			Fvk3a4;
	reg			Fxk3a4;
	reg			Fzk3a4;
	reg			F1l3a4;
	reg			F3l3a4;
	reg			F5l3a4;
	reg			F7l3a4;
	reg			E9l3a4;
	reg			Dbl3a4;
	reg			Cdl3a4;
	reg			Cfl3a4;
	reg			Bhl3a4;
	reg			Ajl3a4;
	reg			Zkl3a4;
	reg			Yml3a4;
	reg			Xol3a4;
	reg			Xql3a4;
	reg			Xsl3a4;
	reg			Xul3a4;
	reg			Xwl3a4;
	reg			Xyl3a4;
	reg			X0m3a4;
	reg			X2m3a4;
	reg			X4m3a4;
	reg			X6m3a4;
	reg			X8m3a4;
	reg			Xam3a4;
	reg			Xcm3a4;
	reg			Xem3a4;
	reg			Xgm3a4;
	reg			Xim3a4;
	reg			Xkm3a4;
	reg			Xmm3a4;
	reg			Xom3a4;
	reg			Xqm3a4;
	reg			Xsm3a4;
	reg			Xum3a4;
	reg			Xwm3a4;
	reg			Xym3a4;
	reg			X0n3a4;
	reg			X2n3a4;
	reg			X4n3a4;
	reg			W6n3a4;
	reg			V8n3a4;
	reg			Uan3a4;
	reg			Tcn3a4;
	reg			Sen3a4;
	reg			Sgn3a4;
	reg			Rin3a4;
	reg			Qkn3a4;
	reg			Pmn3a4;
	reg			Oon3a4;
	reg			Nqn3a4;
	reg			Msn3a4;
	reg			Mun3a4;
	reg			Lwn3a4;
	reg			Kyn3a4;
	reg			J0o3a4;
	reg			I2o3a4;
	reg			H4o3a4;
	reg			H6o3a4;
	reg			H8o3a4;
	reg			Hao3a4;
	reg			Hco3a4;
	reg			Heo3a4;
	reg			Hgo3a4;
	reg			Hio3a4;
	reg			Hko3a4;
	reg			Hmo3a4;
	reg			Hoo3a4;
	reg			Hqo3a4;
	reg			Hso3a4;
	reg			Huo3a4;
	reg			Hwo3a4;
	reg			Hyo3a4;
	reg			H0p3a4;
	reg			H2p3a4;
	reg			H4p3a4;
	reg			H6p3a4;
	reg			H8p3a4;
	reg			Hap3a4;
	reg			Hcp3a4;
	reg			Hep3a4;
	reg			Hgp3a4;
	reg			Hip3a4;
	reg			Hkp3a4;
	reg			Gmp3a4;
	reg			Fop3a4;
	reg			Eqp3a4;
	reg			Dsp3a4;
	reg			Cup3a4;
	reg			Cwp3a4;
	reg			Byp3a4;
	reg			A0q3a4;
	reg			Z1q3a4;
	reg			Y3q3a4;
	reg			X5q3a4;
	reg			W7q3a4;
	reg			W9q3a4;
	reg			Vbq3a4;
	reg			Udq3a4;
	reg			Tfq3a4;
	reg			Shq3a4;
	reg			Rjq3a4;
	reg			Rlq3a4;
	reg			Rnq3a4;
	reg			Rpq3a4;
	reg			Rrq3a4;
	reg			Rtq3a4;
	reg			Rvq3a4;
	reg			Rxq3a4;
	reg			Rzq3a4;
	reg			R1r3a4;
	reg			R3r3a4;
	reg			R5r3a4;
	reg			R7r3a4;
	reg			R9r3a4;
	reg			Qbr3a4;
	reg			Pdr3a4;
	reg			Ofr3a4;
	reg			Ohr3a4;
	reg			Njr3a4;
	reg			Mlr3a4;
	reg			Lnr3a4;
	reg			Kpr3a4;
	reg			Jrr3a4;
	reg			Jtr3a4;
	reg			Jvr3a4;
	reg			Jxr3a4;
	reg			Jzr3a4;
	reg			J1s3a4;
	reg			J3s3a4;
	reg			J5s3a4;
	reg			J7s3a4;
	reg			J9s3a4;
	reg			Jbs3a4;
	reg			Jds3a4;
	reg			Jfs3a4;
	reg			Jhs3a4;
	reg			Jjs3a4;
	reg			Jls3a4;
	reg			Jns3a4;
	reg			Ips3a4;
	reg			Hrs3a4;
	reg			Gts3a4;
	reg			Fvs3a4;
	reg			Exs3a4;
	reg			Dzs3a4;
	reg			C1t3a4;
	reg			C3t3a4;
	reg			C5t3a4;
	reg			C7t3a4;
	reg			C9t3a4;
	reg			Cbt3a4;
	reg			Cdt3a4;
	reg			Cft3a4;
	reg			Cht3a4;
	reg			Cjt3a4;
	reg			Clt3a4;
	reg			Cnt3a4;
	reg			Bpt3a4;
	reg			Art3a4;
	reg			Zst3a4;
	reg			Zut3a4;
	reg			Zwt3a4;
	reg			Yyt3a4;
	reg			X0u3a4;
	reg			W2u3a4;
	reg			V4u3a4;
	reg			U6u3a4;
	reg			T8u3a4;
	reg			Sau3a4;
	reg			Scu3a4;
	reg			Seu3a4;
	reg			Sgu3a4;
	reg			Siu3a4;
	reg			Sku3a4;
	reg			Smu3a4;
	reg			Sou3a4;
	reg			Squ3a4;
	reg			Ssu3a4;
	reg			Suu3a4;
	reg			Swu3a4;
	reg			Syu3a4;
	reg			R0v3a4;
	reg			Q2v3a4;
	reg			P4v3a4;
	reg			P6v3a4;
	reg			O8v3a4;
	reg			Nav3a4;
	reg			Mcv3a4;
	reg			Lev3a4;
	reg			Kgv3a4;
	reg			Kiv3a4;
	reg			Kkv3a4;
	reg			Kmv3a4;
	reg			Kov3a4;
	reg			Kqv3a4;
	reg			Ksv3a4;
	reg			Kuv3a4;
	reg			Kwv3a4;
	reg			Kyv3a4;
	reg			K0w3a4;
	reg			K2w3a4;
	reg			K4w3a4;
	reg			K6w3a4;
	reg			J8w3a4;
	reg			Iaw3a4;
	reg			Hcw3a4;
	reg			Hew3a4;
	reg			Ggw3a4;
	reg			Fiw3a4;
	reg			Ekw3a4;
	reg			Dmw3a4;
	reg			Cow3a4;
	reg			Cqw3a4;
	reg			Csw3a4;
	reg			Cuw3a4;
	reg			Cww3a4;
	reg			Cyw3a4;
	reg			C0x3a4;
	reg			C2x3a4;
	reg			C4x3a4;
	reg			C6x3a4;
	reg			C8x3a4;
	reg			Cax3a4;
	reg			Ccx3a4;
	reg			Cex3a4;
	reg			Bgx3a4;
	reg			Aix3a4;
	reg			Zjx3a4;
	reg			Zlx3a4;
	reg			Ynx3a4;
	reg			Xpx3a4;
	reg			Wrx3a4;
	reg			Vtx3a4;
	reg			Uvx3a4;
	reg			Uxx3a4;
	reg			Uzx3a4;
	reg			U1y3a4;
	reg			U3y3a4;
	reg			U5y3a4;
	reg			U7y3a4;
	reg			U9y3a4;
	reg			Uby3a4;
	reg			Udy3a4;
	reg			Ufy3a4;
	reg			Uhy3a4;
	reg			Ujy3a4;
	reg			Uly3a4;
	reg			Tny3a4;
	reg			Spy3a4;
	reg			Rry3a4;
	reg			Rty3a4;
	reg			Qvy3a4;
	reg			Pxy3a4;
	reg			Ozy3a4;
	reg			N1z3a4;
	reg			M3z3a4;
	reg			M5z3a4;
	reg			M7z3a4;
	reg			M9z3a4;
	reg			Mbz3a4;
	reg			Mdz3a4;
	reg			Mfz3a4;
	reg			Mhz3a4;
	reg			Mjz3a4;
	reg			Mlz3a4;
	reg			Mnz3a4;
	reg			Mpz3a4;
	reg			Mrz3a4;
	reg			Mtz3a4;
	reg			Mvz3a4;
	reg			Mxz3a4;
	reg			Mzz3a4;
	reg			M104a4;
	reg			M304a4;
	reg			M504a4;
	reg			M704a4;
	reg			M904a4;
	reg			Mb04a4;
	reg			Md04a4;
	reg			Mf04a4;
	reg			Mh04a4;
	reg			Mj04a4;
	reg			Ml04a4;
	reg			Mn04a4;
	reg			Mp04a4;
	reg			Mr04a4;
	reg			Lt04a4;
	reg			Kv04a4;
	reg			Kx04a4;
	reg			Kz04a4;
	reg			K114a4;
	reg			K314a4;
	reg			K514a4;
	reg			K714a4;
	reg			K914a4;
	reg			Kb14a4;
	reg			Kd14a4;
	reg			Kf14a4;
	reg			Jh14a4;
	reg			Ij14a4;
	reg			Hl14a4;
	reg			Gn14a4;
	reg			Gp14a4;
	reg			Gr14a4;
	reg			Gt14a4;
	reg			Gv14a4;
	reg			Gx14a4;
	reg			Gz14a4;
	reg			G124a4;
	reg			G324a4;
	reg			G524a4;
	reg			G724a4;
	reg			G924a4;
	reg			Gb24a4;
	reg			Gd24a4;
	reg			Gf24a4;
	reg			Eiwla4;
	reg			Ekwla4;
	reg			Emwla4;
	reg			Dowla4;
	reg			Cqwla4;
	reg			Dswla4;
	reg			Cuwla4;
	reg			Bwwla4;
	reg			Aywla4;
	reg			Zzwla4;
	reg			Z1xla4;
	reg			Z3xla4;
	reg			Z5xla4;
	reg			Z7xla4;
	reg			Z9xla4;
	reg			Zbxla4;
	reg			Zdxla4;
	reg			Zfxla4;
	reg			Zhxla4;
	reg			Zjxla4;
	reg			Zlxla4;
	reg			Znxla4;
	reg			Zpxla4;
	reg			Zrxla4;
	reg			Ztxla4;
	reg			Zvxla4;
	reg			Yxxla4;
	reg			Yzxla4;
	reg			Y1yla4;
	reg			Y3yla4;
	reg			Y5yla4;
	reg			Y7yla4;
	reg			Y9yla4;
	reg			Ybyla4;
	reg			Ydyla4;
	reg			Yfyla4;
	reg			Yhyla4;
	reg			Yjyla4;
	reg			Ylyla4;
	reg			Ynyla4;
	reg			Ypyla4;
	reg			Yryla4;
	reg			Ytyla4;
	reg			Xvyla4;
	reg			Xxyla4;
	reg			Xzyla4;
	reg			X1zla4;
	reg			X3zla4;
	reg			X5zla4;
	reg			X7zla4;
	reg			X9zla4;
	reg			Xbzla4;
	reg			Xdzla4;
	reg			Xfzla4;
	reg			Xhzla4;
	reg			Xjzla4;
	reg			Xlzla4;
	reg			Xnzla4;
	reg			Xpzla4;
	reg			Xrzla4;
	reg			Wtzla4;
	reg			Vvzla4;
	reg			Uxzla4;
	reg			Vzzla4;
	reg			W10ma4;
	reg			T30ma4;
	reg			T50ma4;
	reg			T70ma4;
	reg			T90ma4;
	reg			Tb0ma4;
	reg			Td0ma4;
	reg			Tf0ma4;
	reg			Th0ma4;
	reg			Tj0ma4;
	reg			Tl0ma4;
	reg			Tn0ma4;
	reg			Tp0ma4;
	reg			Tr0ma4;
	reg			Tt0ma4;
	reg			Tv0ma4;
	reg			Tx0ma4;
	reg			Tz0ma4;
	reg			T11ma4;
	reg			Q31ma4;
	reg			Q51ma4;
	reg			Q71ma4;
	reg			Q91ma4;
	reg			Qb1ma4;
	reg			Qd1ma4;
	reg			Qf1ma4;
	reg			Qh1ma4;
	reg			Qj1ma4;
	reg			Ql1ma4;
	reg			Qn1ma4;
	reg			Qp1ma4;
	reg			Qr1ma4;
	reg			Qt1ma4;
	reg			Qv1ma4;
	reg			Qx1ma4;
	reg			Qz1ma4;
	reg			Q12ma4;
	reg			M32ma4;
	reg			L52ma4;
	reg			K72ma4;
	reg			J92ma4;
	reg			Ib2ma4;
	reg			Hd2ma4;
	reg			Gf2ma4;
	reg			Fh2ma4;
	reg			Ej2ma4;
	reg			Dl2ma4;
	reg			Cn2ma4;
	reg			Bp2ma4;
	reg			Ar2ma4;
	reg			Zs2ma4;
	reg			Yu2ma4;
	reg			Xw2ma4;
	reg			Wy2ma4;
	reg			V03ma4;
	reg			U23ma4;
	reg			T43ma4;
	reg			S63ma4;
	reg			R83ma4;
	reg			Qa3ma4;
	reg			Pc3ma4;
	reg			Oe3ma4;
	reg			Ng3ma4;
	reg			Mi3ma4;
	reg			Lk3ma4;
	reg			Km3ma4;
	reg			Jo3ma4;
	reg			Iq3ma4;
	reg			Hs3ma4;
	reg			Gu3ma4;
	reg			Fw3ma4;
	reg			Cy3ma4;
	reg			D04ma4;
	reg			E24ma4;
	reg			F44ma4;
	reg			E64ma4;
	reg			D84ma4;
	reg			Fa4ma4;
	reg			Hc4ma4;
	reg			Je4ma4;
	reg			Lg4ma4;
	reg			Ni4ma4;
	reg			Pk4ma4;
	reg			Qm4ma4;
	reg			Ro4ma4;
	reg			Sq4ma4;
	reg			Ss4ma4;
	reg			Uu4ma4;
	reg			Ww4ma4;
	reg			Yy4ma4;
	reg			A15ma4;
	reg			A35ma4;
	reg			A55ma4;
	reg			A75ma4;
	reg			A95ma4;
	reg			Cb5ma4;
	reg			Ed5ma4;
	reg			Ff5ma4;
	reg			Gh5ma4;
	reg			Hj5ma4;
	reg			Il5ma4;
	reg			Jn5ma4;
	reg			Kp5ma4;
	reg			Lr5ma4;
	reg			Mt5ma4;
	reg			Nv5ma4;
	reg			Ox5ma4;
	reg			Pz5ma4;
	reg			Q16ma4;
	reg			R36ma4;
	reg			S56ma4;
	reg			R76ma4;
	reg			R96ma4;
	reg			Rb6ma4;
	reg			Rd6ma4;
	reg			Rf6ma4;
	reg			Rh6ma4;
	reg			Rj6ma4;
	reg			Rl6ma4;
	reg			Rn6ma4;
	reg			Rp6ma4;
	reg			Rr6ma4;
	reg			Rt6ma4;
	reg			Rv6ma4;
	reg			Rx6ma4;
	reg			Rz6ma4;
	reg			R17ma4;
	reg			R37ma4;
	reg			R57ma4;
	reg			R77ma4;
	reg			T97ma4;
	reg			Vb7ma4;
	reg			Wd7ma4;
	reg			Xf7ma4;
	reg			Zh7ma4;
	reg			Bk7ma4;
	reg			Dm7ma4;
	reg			Fo7ma4;
	reg			Gq7ma4;
	reg			Hs7ma4;
	reg			Iu7ma4;
	reg			Hw7ma4;
	reg			Jy7ma4;
	reg			L08ma4;
	reg			M28ma4;
	reg			O48ma4;
	reg			P68ma4;
	reg			R88ma4;
	reg			Ta8ma4;
	reg			Uc8ma4;
	reg			Ve8ma4;
	wire	[33:0]		Xg8ma4;
	wire	[33:0]		Yi8ma4;

	assign HPROT[1] = 1'b1;
	assign HBURST[2] = 1'b0;
	assign HBURST[1] = 1'b0;
	assign HBURST[0] = 1'b0;
	assign HMASTLOCK = 1'b0;
	assign HSIZE[2] = 1'b0;
	assign HTRANS[0] = 1'b0;
	assign Q34x84 = Db73a4;
	assign Hj5w84 = Ed73a4;
	assign Jd9w84 = Cf73a4;
	assign Js3x84 = Bh73a4;
	assign Aq4w84 = Aj73a4;
	assign Gz4w84 = Yk73a4;
	assign Iv6w84 = Um73a4;
	assign O75w84 = Xo73a4;
	assign Exjw84 = Wq73a4;
	assign Eo5w84 = Ws73a4;
	assign Ol2x84 = Qu73a4;
	assign Th5w84 = Lw73a4;
	assign Geaw84 = Fy73a4;
	assign K6kw84 = F083a4;
	assign Y7xw84 = F283a4;
	assign Nj63a4[4] = F483a4;
	assign I49w84 = B683a4;
	assign Mwiw84 = A883a4;
	assign Ayvw84 = Z983a4;
	assign Tk63a4[25] = Yb83a4;
	assign S8aw84 = Vd83a4;
	assign W0kw84 = Vf83a4;
	assign Sfvw84 = Vh83a4;
	assign O4kw84 = Vj83a4;
	assign C6xw84 = Vl83a4;
	assign Td3x84 = Vn83a4;
	assign Yk0x84 = Sp83a4;
	assign Nj63a4[0] = Rr83a4;
	assign Ke63a4 = Nt83a4;
	assign La3x84 = Kv83a4;
	assign Tm0x84 = Hx83a4;
	assign Ct5w84 = Gz83a4;
	assign Xw6w84 = F193a4;
	assign Oo0x84 = I393a4;
	assign Uu5w84 = H593a4;
	assign Zo2x84 = G793a4;
	assign Bw2x84 = E993a4;
	assign Vx2x84 = Cb93a4;
	assign Me5w84 = Ad93a4;
	assign Tk63a4[2] = Ve93a4;
	assign N29w84 = Rg93a4;
	assign Ruiw84 = Qi93a4;
	assign Fwvw84 = Pk93a4;
	assign Tk63a4[30] = Om93a4;
	assign Yhaw84 = Lo93a4;
	assign D373a4[1] = Lq93a4;
	assign Ws4w84 = Ms93a4;
	assign SLEEPHOLDACKn = Mu93a4;
	assign Qq8x84 = (!Mu93a4);
	assign Tq2x84 = Nw93a4;
	assign Pz2x84 = Ly93a4;
	assign Bg5w84 = J0a3a4;
	assign Yk5w84 = H2a3a4;
	assign Mdxw84 = D4a3a4;
	assign X473a4[10] = Z5a3a4;
	assign Pu63a4[10] = B8a3a4;
	assign Wsiw84 = Daa3a4;
	assign Kuvw84 = Cca3a4;
	assign Tk63a4[15] = Bea3a4;
	assign Gq9w84 = Yfa3a4;
	assign X473a4[16] = Yha3a4;
	assign Pu63a4[16] = Aka3a4;
	assign Vk3x84 = Cma3a4;
	assign P25w84 = Boa3a4;
	assign Cx8w84 = Upa3a4;
	assign Nr4w84 = Tra3a4;
	assign Tk63a4[19] = Pta3a4;
	assign Qx9w84 = Mva3a4;
	assign X473a4[20] = Mxa3a4;
	assign Pu63a4[20] = Oza3a4;
	assign Tk63a4[11] = Q1b3a4;
	assign Wi9w84 = N3b3a4;
	assign X473a4[12] = N5b3a4;
	assign Pu63a4[12] = P7b3a4;
	assign Upjw84 = R9b3a4;
	assign Q4vw84 = Rbb3a4;
	assign Up5w84 = Rdb3a4;
	assign Cakw84 = Lfb3a4;
	assign G2uw84 = Lhb3a4;
	assign Tk63a4[28] = Ljb3a4;
	assign J13x84 = Ilb3a4;
	assign Ap6w84 = Dnb3a4;
	assign Ogjw84 = Cpb3a4;
	assign Kvuw84 = Crb3a4;
	assign Nz63a4[3] = Ctb3a4;
	assign Tk63a4[14] = Dvb3a4;
	assign Ko9w84 = Axb3a4;
	assign Kijw84 = Azb3a4;
	assign Gxuw84 = A1c3a4;
	assign Tk63a4[10] = A3c3a4;
	assign Ah9w84 = X4c3a4;
	assign X473a4[11] = X6c3a4;
	assign Pu63a4[11] = Z8c3a4;
	assign Pu63a4[23] = Bbc3a4;
	assign X1jw84 = Ddc3a4;
	assign Busw84 = Cfc3a4;
	assign Nz63a4[1] = Bhc3a4;
	assign Jq0x84 = Cjc3a4;
	assign Mw5w84 = Blc3a4;
	assign Fn2x84 = Anc3a4;
	assign My6w84 = Yoc3a4;
	assign Ab5w84 = Brc3a4;
	assign Tk63a4[17] = Atc3a4;
	assign Yt9w84 = Xuc3a4;
	assign X473a4[18] = Xwc3a4;
	assign Pu63a4[18] = Zyc3a4;
	assign Tk63a4[9] = B1d3a4;
	assign Ef9w84 = X2d3a4;
	assign I7jw84 = X4d3a4;
	assign Emuw84 = X6d3a4;
	assign Cw3x84 = X8d3a4;
	assign Briw84 = Yad3a4;
	assign X473a4[17] = Xcd3a4;
	assign Pu63a4[17] = Zed3a4;
	assign Tk63a4[16] = Bhd3a4;
	assign Cs9w84 = Yid3a4;
	assign Gkjw84 = Ykd3a4;
	assign Ulww84 = Ymd3a4;
	assign Tk63a4[29] = Yod3a4;
	assign Cgaw84 = Vqd3a4;
	assign D373a4[0] = Vsd3a4;
	assign Tk63a4[5] = Wud3a4;
	assign Y79w84 = Swd3a4;
	assign Nz63a4[0] = Ryd3a4;
	assign Tk63a4[13] = S0e3a4;
	assign Om9w84 = P2e3a4;
	assign Sejw84 = P4e3a4;
	assign Otuw84 = P6e3a4;
	assign Tk63a4[22] = P8e3a4;
	assign E3aw84 = Mae3a4;
	assign Hw63a4[1] = Mce3a4;
	assign Dj0x84 = Lee3a4;
	assign Uj2x84 = Kge3a4;
	assign Wz5w84 = Iie3a4;
	assign Ns2x84 = Hke3a4;
	assign Hu2x84 = Fme3a4;
	assign Nj63a4[2] = Doe3a4;
	assign Nj63a4[3] = Zpe3a4;
	assign Nj63a4[1] = Vre3a4;
	assign Ju4w84 = Rte3a4;
	assign Om5w84 = Pve3a4;
	assign Kcaw84 = Jxe3a4;
	assign Tc2x84 = Jze3a4;
	assign C92x84 = G1f3a4;
	assign W05w84 = G3f3a4;
	assign H95w84 = G5f3a4;
	assign Hyiw84 = F7f3a4;
	assign Vzvw84 = E9f3a4;
	assign Tk63a4[27] = Dbf3a4;
	assign Tk63a4[26] = Adf3a4;
	assign Oaaw84 = Xef3a4;
	assign S2kw84 = Xgf3a4;
	assign Ohvw84 = Xif3a4;
	assign Tk63a4[21] = Xkf3a4;
	assign I1aw84 = Umf3a4;
	assign Mtjw84 = Uof3a4;
	assign I8vw84 = Uqf3a4;
	assign Nj63a4[5] = Usf3a4;
	assign G33x84 = Quf3a4;
	assign Kf3x84 = Rwf3a4;
	assign D69w84 = Oyf3a4;
	assign C0jw84 = N0g3a4;
	assign Q1ww84 = M2g3a4;
	assign Tk63a4[24] = L4g3a4;
	assign W6aw84 = I6g3a4;
	assign Azjw84 = I8g3a4;
	assign Wdvw84 = Iag3a4;
	assign Gpiw84 = Icg3a4;
	assign In4w84 = Heg3a4;
	assign Lo4w84 = Hgg3a4;
	assign Tt6w84 = Jig3a4;
	assign D53x84 = Ikg3a4;
	assign C45w84 = Hmg3a4;
	assign Nx4w84 = Gog3a4;
	assign Ya2x84 = Dqg3a4;
	assign G72x84 = Csg3a4;
	assign K52x84 = Cug3a4;
	assign O32x84 = Cwg3a4;
	assign S12x84 = Cyg3a4;
	assign Wz1x84 = C0h3a4;
	assign Ay1x84 = C2h3a4;
	assign Fw1x84 = C4h3a4;
	assign Ku1x84 = B6h3a4;
	assign Ps1x84 = A8h3a4;
	assign Uq1x84 = Z9h3a4;
	assign Zo1x84 = Ybh3a4;
	assign En1x84 = Xdh3a4;
	assign Jl1x84 = Wfh3a4;
	assign Oj1x84 = Vhh3a4;
	assign Th1x84 = Ujh3a4;
	assign Yf1x84 = Tlh3a4;
	assign Zg6w84 = Snh3a4;
	assign Tk63a4[0] = Sph3a4;
	assign Tk63a4[6] = Orh3a4;
	assign Tk63a4[8] = Kth3a4;
	assign Tk63a4[4] = Gvh3a4;
	assign V55w84 = Cxh3a4;
	assign Uv4w84 = Yyh3a4;
	assign Tk63a4[3] = V0i3a4;
	assign Tk63a4[23] = R2i3a4;
	assign Ig2x84 = O4i3a4;
	assign Bi2x84 = L6i3a4;
	assign S61x84 = I8i3a4;
	assign Uv0x84 = Iai3a4;
	assign Px0x84 = Hci3a4;
	assign Kz0x84 = Gei3a4;
	assign F11x84 = Fgi3a4;
	assign A31x84 = Eii3a4;
	assign W41x84 = Eki3a4;
	assign O81x84 = Emi3a4;
	assign Ka1x84 = Eoi3a4;
	assign Ce1x84 = Eqi3a4;
	assign Gc1x84 = Esi3a4;
	assign Es0x84 = Eui3a4;
	assign Zt0x84 = Dwi3a4;
	assign Ih0x84 = Cyi3a4;
	assign Ey5w84 = Zzi3a4;
	assign O16w84 = Y1j3a4;
	assign G36w84 = X3j3a4;
	assign Y46w84 = W5j3a4;
	assign Q66w84 = V7j3a4;
	assign I86w84 = U9j3a4;
	assign Ba6w84 = Ubj3a4;
	assign Ub6w84 = Udj3a4;
	assign Cc3x84 = Ufj3a4;
	assign Gf6w84 = Rhj3a4;
	assign Kr5w84 = Rjj3a4;
	assign Nd6w84 = Qlj3a4;
	assign C07w84 = Qnj3a4;
	assign Pq6w84 = Tpj3a4;
	assign Es6w84 = Srj3a4;
	assign Km63a4[1] = Rtj3a4;
	assign Km63a4[2] = Qvj3a4;
	assign Km63a4[3] = Pxj3a4;
	assign Km63a4[0] = Ozj3a4;
	assign Tc5w84 = N1k3a4;
	assign Mf0x84 = M3k3a4;
	assign Gyyw84 = M5k3a4;
	assign R3zw84 = L7k3a4;
	assign B0zw84 = K9k3a4;
	assign M5zw84 = Jbk3a4;
	assign W1zw84 = Idk3a4;
	assign H7zw84 = Hfk3a4;
	assign Sczw84 = Ghk3a4;
	assign Ckzw84 = Fjk3a4;
	assign Ylzw84 = Flk3a4;
	assign Qpzw84 = Fnk3a4;
	assign Evzw84 = Fpk3a4;
	assign Wyzw84 = Frk3a4;
	assign K40x84 = Ftk3a4;
	assign G60x84 = Fvk3a4;
	assign C80x84 = Fxk3a4;
	assign Y90x84 = Fzk3a4;
	assign Ub0x84 = F1l3a4;
	assign Unzw84 = F3l3a4;
	assign O20x84 = F5l3a4;
	assign Ybkw84 = F7l3a4;
	assign Tdkw84 = E9l3a4;
	assign Ofkw84 = Dbl3a4;
	assign Uwlw84 = Cdl3a4;
	assign Zkkw84 = Cfl3a4;
	assign Jhkw84 = Bhl3a4;
	assign Umkw84 = Ajl3a4;
	assign Ejkw84 = Zkl3a4;
	assign Pokw84 = Yml3a4;
	assign Aukw84 = Xol3a4;
	assign K1lw84 = Xql3a4;
	assign G3lw84 = Xsl3a4;
	assign Y6lw84 = Xul3a4;
	assign Mclw84 = Xwl3a4;
	assign Eglw84 = Xyl3a4;
	assign Sllw84 = X0m3a4;
	assign Onlw84 = X2m3a4;
	assign Kplw84 = X4m3a4;
	assign Grlw84 = X6m3a4;
	assign Ctlw84 = X8m3a4;
	assign C5lw84 = Xam3a4;
	assign Wjlw84 = Xcm3a4;
	assign O6nw84 = Xem3a4;
	assign Urmw84 = Xgm3a4;
	assign Ufnw84 = Xim3a4;
	assign Ydnw84 = Xkm3a4;
	assign Ccnw84 = Xmm3a4;
	assign Ganw84 = Xom3a4;
	assign K8nw84 = Xqm3a4;
	assign W2nw84 = Xsm3a4;
	assign Ezmw84 = Xum3a4;
	assign Qtmw84 = Xwm3a4;
	assign Ypmw84 = Xym3a4;
	assign Comw84 = X0n3a4;
	assign Sgmw84 = X2n3a4;
	assign Hbmw84 = X4n3a4;
	assign W5mw84 = W6n3a4;
	assign M9mw84 = V8n3a4;
	assign B4mw84 = Uan3a4;
	assign R7mw84 = Tcn3a4;
	assign Mjnw84 = Sen3a4;
	assign G2mw84 = Sgn3a4;
	assign L0mw84 = Rin3a4;
	assign Qylw84 = Qkn3a4;
	assign Ilnw84 = Pmn3a4;
	assign Dnnw84 = Oon3a4;
	assign Yonw84 = Nqn3a4;
	assign E6pw84 = Msn3a4;
	assign Junw84 = Mun3a4;
	assign Tqnw84 = Lwn3a4;
	assign Ewnw84 = Kyn3a4;
	assign Osnw84 = J0o3a4;
	assign Zxnw84 = I2o3a4;
	assign K3ow84 = H4o3a4;
	assign Uaow84 = H6o3a4;
	assign Qcow84 = H8o3a4;
	assign Igow84 = Hao3a4;
	assign Wlow84 = Hco3a4;
	assign Opow84 = Heo3a4;
	assign Cvow84 = Hgo3a4;
	assign Ywow84 = Hio3a4;
	assign Uyow84 = Hko3a4;
	assign Q0pw84 = Hmo3a4;
	assign M2pw84 = Hoo3a4;
	assign Meow84 = Hqo3a4;
	assign Gtow84 = Hso3a4;
	assign Yfqw84 = Huo3a4;
	assign E1qw84 = Hwo3a4;
	assign Epqw84 = Hyo3a4;
	assign Inqw84 = H0p3a4;
	assign Mlqw84 = H2p3a4;
	assign Qjqw84 = H4p3a4;
	assign Uhqw84 = H6p3a4;
	assign Gcqw84 = H8p3a4;
	assign O8qw84 = Hap3a4;
	assign A3qw84 = Hcp3a4;
	assign Izpw84 = Hep3a4;
	assign Mxpw84 = Hgp3a4;
	assign Cqpw84 = Hip3a4;
	assign Rkpw84 = Hkp3a4;
	assign Gfpw84 = Gmp3a4;
	assign Wipw84 = Fop3a4;
	assign Ldpw84 = Eqp3a4;
	assign Bhpw84 = Dsp3a4;
	assign Wsqw84 = Cup3a4;
	assign Qbpw84 = Cwp3a4;
	assign V9pw84 = Byp3a4;
	assign A8pw84 = A0q3a4;
	assign Suqw84 = Z1q3a4;
	assign Nwqw84 = Y3q3a4;
	assign Iyqw84 = X5q3a4;
	assign Ofsw84 = W7q3a4;
	assign T3rw84 = W9q3a4;
	assign D0rw84 = Vbq3a4;
	assign O5rw84 = Udq3a4;
	assign Y1rw84 = Tfq3a4;
	assign J7rw84 = Shq3a4;
	assign Ucrw84 = Rjq3a4;
	assign Ekrw84 = Rlq3a4;
	assign Amrw84 = Rnq3a4;
	assign Sprw84 = Rpq3a4;
	assign Gvrw84 = Rrq3a4;
	assign Yyrw84 = Rtq3a4;
	assign M4sw84 = Rvq3a4;
	assign I6sw84 = Rxq3a4;
	assign E8sw84 = Rzq3a4;
	assign Aasw84 = R1r3a4;
	assign Wbsw84 = R3r3a4;
	assign Wnrw84 = R5r3a4;
	assign Q2sw84 = R7r3a4;
	assign C4uw84 = R9r3a4;
	assign X5uw84 = Qbr3a4;
	assign S7uw84 = Pdr3a4;
	assign Yovw84 = Ofr3a4;
	assign Dduw84 = Ohr3a4;
	assign N9uw84 = Njr3a4;
	assign Yeuw84 = Mlr3a4;
	assign Ibuw84 = Lnr3a4;
	assign Tguw84 = Kpr3a4;
	assign Czuw84 = Jrr3a4;
	assign Kjvw84 = Jtr3a4;
	assign Glvw84 = Jvr3a4;
	assign Acvw84 = Jxr3a4;
	assign Iptw84 = Jzr3a4;
	assign Oatw84 = J1s3a4;
	assign Oytw84 = J3s3a4;
	assign Swtw84 = J5s3a4;
	assign Wutw84 = J7s3a4;
	assign Attw84 = J9s3a4;
	assign Ertw84 = Jbs3a4;
	assign Qltw84 = Jds3a4;
	assign Yhtw84 = Jfs3a4;
	assign S8tw84 = Jhs3a4;
	assign W6tw84 = Jjs3a4;
	assign Mzsw84 = Jls3a4;
	assign Qosw84 = Jns3a4;
	assign Gssw84 = Ips3a4;
	assign Vmsw84 = Hrs3a4;
	assign Lqsw84 = Gts3a4;
	assign Alsw84 = Fvs3a4;
	assign Fjsw84 = Exs3a4;
	assign Khsw84 = Dzs3a4;
	assign Kctw84 = C1t3a4;
	assign Syww84 = C3t3a4;
	assign Yjww84 = C5t3a4;
	assign G4xw84 = C7t3a4;
	assign K2xw84 = C9t3a4;
	assign O0xw84 = Cbt3a4;
	assign Avww84 = Cdt3a4;
	assign Irww84 = Cft3a4;
	assign Ciww84 = Cht3a4;
	assign Ggww84 = Cjt3a4;
	assign W8ww84 = Clt3a4;
	assign L3ww84 = Cnt3a4;
	assign Uqvw84 = Bpt3a4;
	assign Psvw84 = Art3a4;
	assign Qbxw84 = Zst3a4;
	assign Kwyw84 = Zut3a4;
	assign Efxw84 = Zwt3a4;
	assign Pkxw84 = Yyt3a4;
	assign Zgxw84 = X0u3a4;
	assign Kmxw84 = W2u3a4;
	assign Uixw84 = V4u3a4;
	assign Foxw84 = U6u3a4;
	assign Qtxw84 = T8u3a4;
	assign A1yw84 = Sau3a4;
	assign W2yw84 = Scu3a4;
	assign O6yw84 = Seu3a4;
	assign Ccyw84 = Sgu3a4;
	assign Ufyw84 = Siu3a4;
	assign Ilyw84 = Sku3a4;
	assign Enyw84 = Smu3a4;
	assign Apyw84 = Sou3a4;
	assign Wqyw84 = Squ3a4;
	assign Ssyw84 = Ssu3a4;
	assign S4yw84 = Suu3a4;
	assign Mjyw84 = Swu3a4;
	assign Ujaw84 = Syu3a4;
	assign Plaw84 = R0v3a4;
	assign Knaw84 = Q2v3a4;
	assign Q4cw84 = P4v3a4;
	assign Vsaw84 = P6v3a4;
	assign Fpaw84 = O8v3a4;
	assign Quaw84 = Nav3a4;
	assign Araw84 = Mcv3a4;
	assign Lwaw84 = Lev3a4;
	assign W1bw84 = Kgv3a4;
	assign G9bw84 = Kiv3a4;
	assign Cbbw84 = Kkv3a4;
	assign Uebw84 = Kmv3a4;
	assign Ikbw84 = Kov3a4;
	assign Aobw84 = Kqv3a4;
	assign Otbw84 = Ksv3a4;
	assign Kvbw84 = Kuv3a4;
	assign Gxbw84 = Kwv3a4;
	assign Czbw84 = Kyv3a4;
	assign Y0cw84 = K0w3a4;
	assign Ycbw84 = K2w3a4;
	assign Srbw84 = K4w3a4;
	assign M6cw84 = K6w3a4;
	assign H8cw84 = J8w3a4;
	assign Cacw84 = Iaw3a4;
	assign Irdw84 = Hcw3a4;
	assign Nfcw84 = Hew3a4;
	assign Xbcw84 = Ggw3a4;
	assign Ihcw84 = Fiw3a4;
	assign Sdcw84 = Ekw3a4;
	assign Djcw84 = Dmw3a4;
	assign Oocw84 = Cow3a4;
	assign Yvcw84 = Cqw3a4;
	assign Uxcw84 = Csw3a4;
	assign M1dw84 = Cuw3a4;
	assign A7dw84 = Cww3a4;
	assign Sadw84 = Cyw3a4;
	assign Ggdw84 = C0x3a4;
	assign Cidw84 = C2x3a4;
	assign Yjdw84 = C4x3a4;
	assign Uldw84 = C6x3a4;
	assign Qndw84 = C8x3a4;
	assign Qzcw84 = Cax3a4;
	assign Kedw84 = Ccx3a4;
	assign O2hw84 = Cex3a4;
	assign J4hw84 = Bgx3a4;
	assign E6hw84 = Aix3a4;
	assign Kniw84 = Zjx3a4;
	assign Pbhw84 = Zlx3a4;
	assign Z7hw84 = Ynx3a4;
	assign Kdhw84 = Xpx3a4;
	assign U9hw84 = Wrx3a4;
	assign Ffhw84 = Vtx3a4;
	assign Qkhw84 = Uvx3a4;
	assign Ashw84 = Uxx3a4;
	assign Wthw84 = Uzx3a4;
	assign Oxhw84 = U1y3a4;
	assign C3iw84 = U3y3a4;
	assign U6iw84 = U5y3a4;
	assign Iciw84 = U7y3a4;
	assign Eeiw84 = U9y3a4;
	assign Agiw84 = Uby3a4;
	assign Whiw84 = Udy3a4;
	assign Sjiw84 = Ufy3a4;
	assign Svhw84 = Uhy3a4;
	assign Maiw84 = Ujy3a4;
	assign Wffw84 = Uly3a4;
	assign Rhfw84 = Tny3a4;
	assign Mjfw84 = Spy3a4;
	assign S0hw84 = Rry3a4;
	assign Xofw84 = Rty3a4;
	assign Hlfw84 = Qvy3a4;
	assign Sqfw84 = Pxy3a4;
	assign Cnfw84 = Ozy3a4;
	assign Nsfw84 = N1z3a4;
	assign Yxfw84 = M3z3a4;
	assign I5gw84 = M5z3a4;
	assign E7gw84 = M7z3a4;
	assign Wagw84 = M9z3a4;
	assign Kggw84 = Mbz3a4;
	assign Ckgw84 = Mdz3a4;
	assign Qpgw84 = Mfz3a4;
	assign Mrgw84 = Mhz3a4;
	assign Itgw84 = Mjz3a4;
	assign Evgw84 = Mlz3a4;
	assign Axgw84 = Mnz3a4;
	assign A9gw84 = Mpz3a4;
	assign Ungw84 = Mrz3a4;
	assign C1fw84 = Mtz3a4;
	assign Imew84 = Mvz3a4;
	assign Iafw84 = Mxz3a4;
	assign M8fw84 = Mzz3a4;
	assign Q6fw84 = M104a4;
	assign U4fw84 = M304a4;
	assign Y2fw84 = M504a4;
	assign Kxew84 = M704a4;
	assign Stew84 = M904a4;
	assign Eoew84 = Mb04a4;
	assign Mkew84 = Md04a4;
	assign Qiew84 = Mf04a4;
	assign Cdew84 = Mh04a4;
	assign Saww84 = Mj04a4;
	assign Yrpw84 = Ml04a4;
	assign Oimw84 = Mn04a4;
	assign I1tw84 = Mp04a4;
	assign Mvxw84 = Mr04a4;
	assign Oezw84 = Lt04a4;
	assign S3bw84 = Kv04a4;
	assign Kqcw84 = Kx04a4;
	assign Wvkw84 = Kz04a4;
	assign G5ow84 = K114a4;
	assign Uzfw84 = K314a4;
	assign Mmhw84 = K514a4;
	assign E9jw84 = K714a4;
	assign Qerw84 = K914a4;
	assign Aouw84 = Kb14a4;
	assign Gbew84 = Kd14a4;
	assign K0ew84 = Kf14a4;
	assign A4ew84 = Jh14a4;
	assign Pydw84 = Ij14a4;
	assign F2ew84 = Hl14a4;
	assign Aefw84 = Gn14a4;
	assign Gzew84 = Gp14a4;
	assign Mntw84 = Gr14a4;
	assign S00x84 = Gt14a4;
	assign S4nw84 = Gv14a4;
	assign Ceqw84 = Gx14a4;
	assign Wwww84 = Gz14a4;
	assign Eavw84 = G124a4;
	assign U0sw84 = G324a4;
	assign Krow84 = G524a4;
	assign Ailw84 = G724a4;
	assign Qhyw84 = G924a4;
	assign Wpbw84 = Gb24a4;
	assign Ocdw84 = Gd24a4;
	assign Ylgw84 = Gf24a4;
	assign Q8iw84 = Eiwla4;
	assign Ivjw84 = Ekwla4;
	assign Zudw84 = Emwla4;
	assign Xy8w84 = Dowla4;
	assign Vs63a4[1] = Cqwla4;
	assign Etdw84 = Dswla4;
	assign Uwdw84 = Cuwla4;
	assign S09w84 = Bwwla4;
	assign V5ew84 = Aywla4;
	assign Y0vw84 = Zzwla4;
	assign Orrw84 = Z1xla4;
	assign Cmjw84 = Z3xla4;
	assign Kzhw84 = Z5xla4;
	assign Scgw84 = Z7xla4;
	assign Aqew84 = Z9xla4;
	assign Eiow84 = Zbxla4;
	assign U8lw84 = Zdxla4;
	assign I3dw84 = Zfxla4;
	assign Qgbw84 = Zhxla4;
	assign Mrzw84 = Zjxla4;
	assign K8yw84 = Zlxla4;
	assign Getw84 = Znxla4;
	assign Mvmw84 = Zpxla4;
	assign W4qw84 = Zrxla4;
	assign Qnww84 = Ztxla4;
	assign Hk6w84 = Zvxla4;
	assign Ocww84 = Yxxla4;
	assign Wpuw84 = Yzxla4;
	assign Mgrw84 = Y1yla4;
	assign Abjw84 = Y3yla4;
	assign Iohw84 = Y5yla4;
	assign Q1gw84 = Y7yla4;
	assign Yeew84 = Y9yla4;
	assign Utpw84 = Ybyla4;
	assign C7ow84 = Ydyla4;
	assign Kkmw84 = Yfyla4;
	assign Sxkw84 = Yhyla4;
	assign Gscw84 = Yjyla4;
	assign O5bw84 = Ylyla4;
	assign Kgzw84 = Ynyla4;
	assign Ixxw84 = Ypyla4;
	assign E3tw84 = Yryla4;
	assign Wl6w84 = Ytyla4;
	assign G8kw84 = Xvyla4;
	assign Oliw84 = Xxyla4;
	assign Wygw84 = Xzyla4;
	assign Ecfw84 = X1zla4;
	assign Mpdw84 = X3zla4;
	assign U2cw84 = X5zla4;
	assign Yulw84 = X7zla4;
	assign I4pw84 = X9zla4;
	assign Sdsw84 = Xbzla4;
	assign Cnvw84 = Xdzla4;
	assign U9xw84 = Xfzla4;
	assign Arqw84 = Xhzla4;
	assign Qhnw84 = Xjzla4;
	assign Ouyw84 = Xlzla4;
	assign Qd0x84 = Xnzla4;
	assign K0uw84 = Xpzla4;
	assign Ln6w84 = Xrzla4;
	assign Si6w84 = Wtzla4;
	assign Y63x84 = Vvzla4;
	assign Pu63a4[0] = Uxzla4;
	assign Pu63a4[3] = Vzzla4;
	assign Tk63a4[18] = W10ma4;
	assign Uv9w84 = T30ma4;
	assign U2vw84 = T50ma4;
	assign Ktrw84 = T70ma4;
	assign Ynjw84 = T90ma4;
	assign G1iw84 = Tb0ma4;
	assign Oegw84 = Td0ma4;
	assign Wrew84 = Tf0ma4;
	assign Akow84 = Th0ma4;
	assign Qalw84 = Tj0ma4;
	assign E5dw84 = Tl0ma4;
	assign Mibw84 = Tn0ma4;
	assign Itzw84 = Tp0ma4;
	assign Gayw84 = Tr0ma4;
	assign Cgtw84 = Tt0ma4;
	assign Ixmw84 = Tv0ma4;
	assign S6qw84 = Tx0ma4;
	assign Mpww84 = Tz0ma4;
	assign Tk63a4[12] = T11ma4;
	assign Sk9w84 = Q31ma4;
	assign Keww84 = Q51ma4;
	assign Qvpw84 = Q71ma4;
	assign Gmmw84 = Q91ma4;
	assign A5tw84 = Qb1ma4;
	assign Ezxw84 = Qd1ma4;
	assign Gizw84 = Qf1ma4;
	assign K7bw84 = Qh1ma4;
	assign Cucw84 = Qj1ma4;
	assign Ozkw84 = Ql1ma4;
	assign Y8ow84 = Qn1ma4;
	assign Ugew84 = Qp1ma4;
	assign M3gw84 = Qr1ma4;
	assign Eqhw84 = Qt1ma4;
	assign Wcjw84 = Qv1ma4;
	assign Iirw84 = Qx1ma4;
	assign Sruw84 = Qz1ma4;
	assign Tk63a4[7] = Q12ma4;
	assign Ob9w84 = M32ma4;
	assign B7ww84 = L52ma4;
	assign Jkuw84 = K72ma4;
	assign Zarw84 = J92ma4;
	assign N5jw84 = Ib2ma4;
	assign Vihw84 = Hd2ma4;
	assign Dwfw84 = Gf2ma4;
	assign L9ew84 = Fh2ma4;
	assign Hopw84 = Ej2ma4;
	assign P1ow84 = Dl2ma4;
	assign Xemw84 = Cn2ma4;
	assign Fskw84 = Bp2ma4;
	assign Tmcw84 = Ar2ma4;
	assign B0bw84 = Zs2ma4;
	assign Xazw84 = Yu2ma4;
	assign Vrxw84 = Xw2ma4;
	assign Rxsw84 = Wy2ma4;
	assign Oiuw84 = V03ma4;
	assign E9rw84 = U23ma4;
	assign S3jw84 = T43ma4;
	assign Ahhw84 = S63ma4;
	assign Iufw84 = R83ma4;
	assign Q7ew84 = Qa3ma4;
	assign Uznw84 = Pc3ma4;
	assign Kqkw84 = Oe3ma4;
	assign Ykcw84 = Ng3ma4;
	assign Gyaw84 = Mi3ma4;
	assign C9zw84 = Lk3ma4;
	assign Aqxw84 = Km3ma4;
	assign Wvsw84 = Jo3ma4;
	assign Cdmw84 = Iq3ma4;
	assign Mmpw84 = Hs3ma4;
	assign G5ww84 = Gu3ma4;
	assign Tk63a4[20] = Fw3ma4;
	assign Wz3x84 = Cy3ma4;
	assign Zx3x84 = D04ma4;
	assign T14x84 = E24ma4;
	assign Xx63a4[0] = F44ma4;
	assign Xx63a4[1] = E64ma4;
	assign N54x84 = (!D84ma4);
	assign Eu3x84 = Fa4ma4;
	assign S54x84 = (!Hc4ma4);
	assign X54x84 = (!Je4ma4);
	assign Oo3x84 = Lg4ma4;
	assign Qm3x84 = Ni4ma4;
	assign Mq3x84 = Pk4ma4;
	assign Nz63a4[6] = Qm4ma4;
	assign Nz63a4[7] = Ro4ma4;
	assign R83x84 = Sq4ma4;
	assign K873a4[1] = Ss4ma4;
	assign K873a4[0] = Uu4ma4;
	assign K873a4[2] = Ww4ma4;
	assign K873a4[3] = Yy4ma4;
	assign R673a4[1] = A15ma4;
	assign R673a4[2] = A35ma4;
	assign R673a4[3] = A55ma4;
	assign R673a4[0] = A75ma4;
	assign X473a4[15] = A95ma4;
	assign Pu63a4[15] = Cb5ma4;
	assign X473a4[9] = Ed5ma4;
	assign Pu63a4[9] = Ff5ma4;
	assign X473a4[7] = Gh5ma4;
	assign Pu63a4[7] = Hj5ma4;
	assign X473a4[6] = Il5ma4;
	assign Pu63a4[6] = Jn5ma4;
	assign X473a4[5] = Kp5ma4;
	assign Pu63a4[5] = Lr5ma4;
	assign X473a4[4] = Mt5ma4;
	assign Pu63a4[4] = Nv5ma4;
	assign X473a4[3] = Ox5ma4;
	assign X473a4[2] = Pz5ma4;
	assign X473a4[1] = Q16ma4;
	assign X473a4[0] = R36ma4;
	assign T99w84 = S56ma4;
	assign A5aw84 = R76ma4;
	assign Mz9w84 = R96ma4;
	assign Etww84 = Rb6ma4;
	assign Kaqw84 = Rd6ma4;
	assign A1nw84 = Rf6ma4;
	assign Ujtw84 = Rh6ma4;
	assign Ydyw84 = Rj6ma4;
	assign Axzw84 = Rl6ma4;
	assign Embw84 = Rn6ma4;
	assign W8dw84 = Rp6ma4;
	assign Ielw84 = Rr6ma4;
	assign Snow84 = Rt6ma4;
	assign Ovew84 = Rv6ma4;
	assign Gigw84 = Rx6ma4;
	assign Y4iw84 = Rz6ma4;
	assign Qrjw84 = R17ma4;
	assign Cxrw84 = R37ma4;
	assign M6vw84 = R57ma4;
	assign X473a4[21] = R77ma4;
	assign Pu63a4[21] = T97ma4;
	assign X473a4[8] = Vb7ma4;
	assign Pu63a4[8] = Wd7ma4;
	assign X473a4[13] = Xf7ma4;
	assign Pu63a4[13] = Zh7ma4;
	assign X473a4[19] = Bk7ma4;
	assign Pu63a4[19] = Dm7ma4;
	assign Pu63a4[2] = Fo7ma4;
	assign Pu63a4[1] = Gq7ma4;
	assign Vs63a4[0] = Hs7ma4;
	assign Hw63a4[0] = Iu7ma4;
	assign X473a4[22] = Hw7ma4;
	assign Pu63a4[22] = Jy7ma4;
	assign Nz63a4[4] = L08ma4;
	assign X473a4[23] = M28ma4;
	assign Nz63a4[5] = O48ma4;
	assign X473a4[14] = P68ma4;
	assign Pu63a4[14] = R88ma4;
	assign Nz63a4[2] = Ta8ma4;
	assign Bh3x84 = Uc8ma4;
	assign SYSRESETREQ = Ve8ma4;
	assign C64x84 = (!Ve8ma4);
	assign H173a4 = (Pu63a4 - 1);
	assign Cr63a4 = ({Tk63a4[30:2], V55w84, Tk63a4[0]} + 1);
	assign {Ao63a4, Fa73a4} = ({Tk63a4[30:2], Me2x84} + 1);
	assign Xg8ma4 = ({{E29x84, S39x84, G59x84, U69x84, I89x84, W99x84,
		Xc9x84, Le9x84, Zf9x84, Nh9x84, Bj9x84, Pk9x84, Dm9x84, Rn9x84,
		Fp9x84, Tq9x84, Hs9x84, Vt9x84, Jv9x84, Xw9x84, Ly9x84, Zz9x84,
		N1ax84, B3ax84, P4ax84, D6ax84, Et8x84, Ru8x84, Ew8x84, Rx8x84,
		Ez8x84, R09x84, Kb9x84}, 1'b0} + {{1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
		1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
		1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
		1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, G37w84}, 1'b1});
	assign {S17w84, Qp63a4} = Xg8ma4[33:1];
	assign Yi8ma4 = ({{1'b0, Gv8w84, Kt8w84, Or8w84, Sp8w84, Wn8w84, Am8w84,
		Ek8w84, Ii8w84, Mg8w84, Qe8w84, Uc8w84, Ya8w84, C98w84, G78w84,
		K58w84, O38w84, S18w84, Wz7w84, Ay7w84, Ew7w84, Iu7w84, Ms7w84,
		Rq7w84, Wo7w84, Bn7w84, Gl7w84, Lj7w84, Qh7w84, Vf7w84, Ae7w84,
		Fc7w84, Ka7w84}, 1'b0} + {{1'b0, Gqax84, H9ax84, A9ax84, V9ax84,
		Hg63a4, O87w84, Ag63a4, O9ax84, Qh63a4, Jh63a4, Vg63a4, Og63a4,
		Qaax84, Xaax84, Caax84, Ch63a4, Si63a4, Li63a4, Ei63a4, Jaax84,
		Zi63a4, Xh63a4, R7ax84, T8ax84, Gj63a4, M8ax84, F8ax84, Y7ax84,
		Ys8x84, Tf63a4, T67w84, Y47w84}, 1'b1});
	assign {E29x84, S39x84, G59x84, U69x84, I89x84, W99x84, Xc9x84, Le9x84, 
		Zf9x84, Nh9x84, Bj9x84, Pk9x84, Dm9x84, Rn9x84, Fp9x84, Tq9x84, 
		Hs9x84, Vt9x84, Jv9x84, Xw9x84, Ly9x84, Zz9x84, N1ax84, B3ax84, 
		P4ax84, D6ax84, Et8x84, Ru8x84, Ew8x84, Rx8x84, Ez8x84, R09x84, 
		Kb9x84} = Yi8ma4[33:1];
	assign Me2x84 = (~(Uqax84 & Brax84));
	assign Brax84 = (~(Irax84 & Tk63a4[0]));
	assign Irax84 = (Prax84 & Wrax84);
	assign Uqax84 = (~(Dsax84 & V55w84));
	assign Rq7w84 = (~(Ksax84 | Rsax84));
	assign Wo7w84 = (~(Ysax84 | Ksax84));
	assign Bn7w84 = (~(Ftax84 | Ksax84));
	assign Gl7w84 = (~(Mtax84 | Ksax84));
	assign Lj7w84 = (~(Ttax84 | Ksax84));
	assign Qh7w84 = (~(Auax84 | Ksax84));
	assign Vf7w84 = (~(Huax84 | Ksax84));
	assign Kt8w84 = (~(Ouax84 | Ksax84));
	assign Ae7w84 = (Vuax84 & Cvax84);
	assign Cvax84 = (~(Jvax84 & Qvax84));
	assign Jvax84 = (~(Xvax84 | Ewax84));
	assign Vuax84 = (~(Lwax84 | Ksax84));
	assign Or8w84 = (~(Swax84 | Ksax84));
	assign Sp8w84 = (~(Zwax84 | Ksax84));
	assign Wn8w84 = (~(Gxax84 | Ksax84));
	assign Am8w84 = (~(Nxax84 | Ksax84));
	assign Ek8w84 = (~(Uxax84 | Ksax84));
	assign Ii8w84 = (~(Byax84 | Ksax84));
	assign Mg8w84 = (~(Iyax84 | Ksax84));
	assign Qe8w84 = (~(Pyax84 | Ksax84));
	assign Uc8w84 = (~(Wyax84 | Ksax84));
	assign Ya8w84 = (~(Dzax84 | Ksax84));
	assign Fc7w84 = (~(Kzax84 | Ksax84));
	assign C98w84 = (~(Rzax84 | Ksax84));
	assign G78w84 = (~(Yzax84 | Ksax84));
	assign K58w84 = (~(F0bx84 | Ksax84));
	assign O38w84 = (~(M0bx84 | Ksax84));
	assign S18w84 = (~(T0bx84 | Ksax84));
	assign Wz7w84 = (~(A1bx84 | Ksax84));
	assign Ay7w84 = (~(H1bx84 | Ksax84));
	assign Ew7w84 = (~(O1bx84 | Ksax84));
	assign Iu7w84 = (~(V1bx84 | Ksax84));
	assign Ms7w84 = (~(C2bx84 | Ksax84));
	assign Ka7w84 = (~(J2bx84 | Ksax84));
	assign Ksax84 = (!Q2bx84);
	assign G37w84 = (~(X2bx84 & E3bx84));
	assign E3bx84 = (~(L3bx84 & S3bx84));
	assign S3bx84 = (Z3bx84 & G4bx84);
	assign Z3bx84 = (~(N4bx84 & U4bx84));
	assign U4bx84 = (B5bx84 | Zo2x84);
	assign L3bx84 = (Th5w84 & I5bx84);
	assign X2bx84 = (~(Ol2x84 & P5bx84));
	assign P5bx84 = (~(W5bx84 & D6bx84));
	assign D6bx84 = (K6bx84 & R6bx84);
	assign R6bx84 = (~(Y6bx84 & F7bx84));
	assign K6bx84 = (M7bx84 & T7bx84);
	assign M7bx84 = (~(A8bx84 & H8bx84));
	assign H8bx84 = (~(B5bx84 | G4bx84));
	assign A8bx84 = (~(N4bx84 | O8bx84));
	assign W5bx84 = (V8bx84 & C9bx84);
	assign C9bx84 = (J9bx84 | Ewax84);
	assign Ss8x84 = (~(Q9bx84 & X9bx84));
	assign X9bx84 = (~(Eabx84 & Labx84));
	assign Labx84 = (~(Sabx84 & Zabx84));
	assign Zabx84 = (Gbbx84 & Nbbx84);
	assign Nbbx84 = (~(Mw5w84 & Ubbx84));
	assign Ubbx84 = (~(Bcbx84 & Icbx84));
	assign Icbx84 = (~(Pcbx84 & Wcbx84));
	assign Gbbx84 = (~(Ba6w84 & Ddbx84));
	assign Ddbx84 = (~(Kdbx84 & Rdbx84));
	assign Sabx84 = (Ydbx84 & Febx84);
	assign Febx84 = (Mebx84 | Tebx84);
	assign Q9bx84 = (~(C07w84 & Afbx84));
	assign Afbx84 = (~(Eabx84 & Hfbx84));
	assign Hfbx84 = (~(Ofbx84 & Vfbx84));
	assign Ms8x84 = (~(Cgbx84 & Jgbx84));
	assign Jgbx84 = (~(My6w84 & Qgbx84));
	assign Qgbx84 = (~(Xgbx84 & Ehbx84));
	assign Ehbx84 = (~(Xw6w84 & Ofbx84));
	assign Cgbx84 = (~(Eabx84 & Lhbx84));
	assign Lhbx84 = (~(Shbx84 & Zhbx84));
	assign Zhbx84 = (Gibx84 & Nibx84);
	assign Nibx84 = (~(Uu5w84 & Uibx84));
	assign Gibx84 = (Bjbx84 & Rdbx84);
	assign Bjbx84 = (Tebx84 | Ijbx84);
	assign Shbx84 = (Ydbx84 & Pjbx84);
	assign Pjbx84 = (Mebx84 | Wcbx84);
	assign Gs8x84 = (~(Wjbx84 & Dkbx84));
	assign Dkbx84 = (Kkbx84 | Xgbx84);
	assign Xgbx84 = (Eabx84 & Rkbx84);
	assign Rkbx84 = (~(Iv6w84 & Ofbx84));
	assign Ofbx84 = (~(Ykbx84 & Flbx84));
	assign Flbx84 = (~(Mlbx84 & Fn2x84));
	assign Ykbx84 = (Tlbx84 & Ambx84);
	assign Wjbx84 = (~(Eabx84 & Hmbx84));
	assign Hmbx84 = (~(Ombx84 & Vmbx84));
	assign Vmbx84 = (Cnbx84 & Jnbx84);
	assign Jnbx84 = (~(Ct5w84 & Uibx84));
	assign Cnbx84 = (Qnbx84 & Rdbx84);
	assign Qnbx84 = (Wcbx84 | Ijbx84);
	assign Ombx84 = (Ydbx84 & Xnbx84);
	assign Xnbx84 = (Eobx84 | Mebx84);
	assign As8x84 = (Lobx84 | Sobx84);
	assign Sobx84 = (Zobx84 & Gpbx84);
	assign Zobx84 = (~(Npbx84 & Upbx84));
	assign Upbx84 = (~(Bqbx84 & Iqbx84));
	assign Bqbx84 = (~(Pqbx84 | Wqbx84));
	assign Npbx84 = (~(Drbx84 & Krbx84));
	assign Krbx84 = (~(Zo2x84 & Rrbx84));
	assign Rrbx84 = (Yrbx84 | Bw2x84);
	assign Lobx84 = (HREADY ? Fsbx84 : Pz2x84);
	assign Fsbx84 = (~(Msbx84 & Tsbx84));
	assign Tsbx84 = (Atbx84 & Htbx84);
	assign Htbx84 = (Otbx84 & Vtbx84);
	assign Vtbx84 = (Cubx84 & Jubx84);
	assign Otbx84 = (Qubx84 & Xubx84);
	assign Qubx84 = (~(Evbx84 & Lvbx84));
	assign Lvbx84 = (~(Svbx84 & Zvbx84));
	assign Zvbx84 = (~(Gwbx84 & Q66w84));
	assign Svbx84 = (Ba6w84 | Gf6w84);
	assign Atbx84 = (Nwbx84 & Uwbx84);
	assign Uwbx84 = (Bxbx84 & Ixbx84);
	assign Ixbx84 = (~(Pxbx84 & Wxbx84));
	assign Wxbx84 = (~(Dybx84 & Kybx84));
	assign Kybx84 = (Rybx84 | Yybx84);
	assign Bxbx84 = (~(Tq2x84 & Fzbx84));
	assign Fzbx84 = (~(Mzbx84 & Tzbx84));
	assign Tzbx84 = (A0cx84 | Yybx84);
	assign Nwbx84 = (H0cx84 & O0cx84);
	assign O0cx84 = (~(Gf6w84 & V0cx84));
	assign V0cx84 = (~(C1cx84 & J1cx84));
	assign J1cx84 = (Q1cx84 | Gpbx84);
	assign C1cx84 = (X1cx84 & E2cx84);
	assign X1cx84 = (~(L2cx84 & S2cx84));
	assign S2cx84 = (~(Z2cx84 & G3cx84));
	assign G3cx84 = (N3cx84 | Eobx84);
	assign Z2cx84 = (~(U3cx84 & B4cx84));
	assign H0cx84 = (I4cx84 | E2cx84);
	assign Msbx84 = (P4cx84 & W4cx84);
	assign W4cx84 = (D5cx84 & K5cx84);
	assign K5cx84 = (R5cx84 & Y5cx84);
	assign Y5cx84 = (F6cx84 | Nd6w84);
	assign D5cx84 = (M6cx84 & T6cx84);
	assign T6cx84 = (~(A7cx84 & Wqbx84));
	assign P4cx84 = (H7cx84 & O7cx84);
	assign O7cx84 = (Gz4w84 ? C8cx84 : V7cx84);
	assign C8cx84 = (J8cx84 & Q8cx84);
	assign Q8cx84 = (~(X8cx84 & E9cx84));
	assign V7cx84 = (L9cx84 & S9cx84);
	assign S9cx84 = (Z9cx84 & Gacx84);
	assign Gacx84 = (~(Nacx84 & Uacx84));
	assign Z9cx84 = (Bbcx84 & B5bx84);
	assign Bbcx84 = (Rybx84 | Tq2x84);
	assign L9cx84 = (Ibcx84 & Pbcx84);
	assign Pbcx84 = (Wbcx84 | Ewax84);
	assign H7cx84 = (Dccx84 & Kccx84);
	assign Kccx84 = (Ambx84 | Ewax84);
	assign Ur8x84 = (~(Rccx84 & Yccx84));
	assign Yccx84 = (~(Fdcx84 & Mdcx84));
	assign Mdcx84 = (~(Tdcx84 & Aecx84));
	assign Aecx84 = (~(G36w84 & Hecx84));
	assign Hecx84 = (~(Oecx84 & Vecx84));
	assign Vecx84 = (Cfcx84 | Tebx84);
	assign Tdcx84 = (Jfcx84 | Qfcx84);
	assign Rccx84 = (~(Tt6w84 & Xfcx84));
	assign Xfcx84 = (~(Fdcx84 & Egcx84));
	assign Egcx84 = (~(Lgcx84 & Sgcx84));
	assign Or8x84 = (~(Zgcx84 & Ghcx84));
	assign Ghcx84 = (~(Fdcx84 & Nhcx84));
	assign Nhcx84 = (~(Uhcx84 & Bicx84));
	assign Bicx84 = (Iicx84 | Qfcx84);
	assign Uhcx84 = (~(O16w84 & Picx84));
	assign Zgcx84 = (~(Es6w84 & Wicx84));
	assign Wicx84 = (~(Fdcx84 & Djcx84));
	assign Djcx84 = (~(Lgcx84 & Kjcx84));
	assign Ir8x84 = (~(Rjcx84 & Yjcx84));
	assign Yjcx84 = (~(Pq6w84 & Fkcx84));
	assign Fkcx84 = (~(Fdcx84 & Mkcx84));
	assign Mkcx84 = (~(Lgcx84 & Tkcx84));
	assign Rjcx84 = (~(Fdcx84 & Alcx84));
	assign Alcx84 = (~(Hlcx84 & Olcx84));
	assign Olcx84 = (Vlcx84 & Cmcx84);
	assign Cmcx84 = (Jmcx84 | Qfcx84);
	assign Vlcx84 = (~(Wz5w84 & Picx84));
	assign Hlcx84 = (Qmcx84 & Xmcx84);
	assign Xmcx84 = (~(Zt0x84 & Encx84));
	assign Qmcx84 = (Lncx84 | Tebx84);
	assign Cr8x84 = (Sncx84 | Zncx84);
	assign Zncx84 = (Gocx84 & Nocx84);
	assign Gocx84 = (~(Uocx84 | Bpcx84));
	assign Sncx84 = (Ppcx84 ? Ipcx84 : Hj5w84);
	assign Ppcx84 = (~(Wpcx84 | Uocx84));
	assign Uocx84 = (Dqcx84 & Kqcx84);
	assign Kqcx84 = (~(Rqcx84 & Qvax84));
	assign Rqcx84 = (~(Yqcx84 | Ewax84));
	assign Dqcx84 = (~(Frcx84 & Mrcx84));
	assign Ipcx84 = (Trcx84 & Ascx84);
	assign Trcx84 = (!Hscx84);
	assign Wq8x84 = (Oscx84 | Vscx84);
	assign Vscx84 = (Ctcx84 & Jtcx84);
	assign Ctcx84 = (~(Qtcx84 | Xtcx84));
	assign Oscx84 = (HREADY ? Eucx84 : Gz4w84);
	assign Eucx84 = (~(Lucx84 & Sucx84));
	assign Sucx84 = (Zucx84 & Gvcx84);
	assign Gvcx84 = (~(Mlbx84 & Nvcx84));
	assign Nvcx84 = (~(Uvcx84 & Bwcx84));
	assign Bwcx84 = (~(Bw2x84 & Iwcx84));
	assign Iwcx84 = (~(Pwcx84 & Wwcx84));
	assign Wwcx84 = (~(Fn2x84 & Dxcx84));
	assign Dxcx84 = (~(Kxcx84 & Rxcx84));
	assign Rxcx84 = (Yxcx84 | Fycx84);
	assign Pwcx84 = (Mycx84 | Fycx84);
	assign Uvcx84 = (Tycx84 & Azcx84);
	assign Azcx84 = (~(Hzcx84 & Ozcx84));
	assign Hzcx84 = (~(Vzcx84 | Ewax84));
	assign Tycx84 = (~(C0dx84 & J0dx84));
	assign Zucx84 = (Q0dx84 & X0dx84);
	assign X0dx84 = (~(E1dx84 & L1dx84));
	assign L1dx84 = (~(S1dx84 & Z1dx84));
	assign Z1dx84 = (~(G2dx84 & N2dx84));
	assign N2dx84 = (U2dx84 & Ln6w84);
	assign U2dx84 = (~(B3dx84 | Ewax84));
	assign G2dx84 = (I3dx84 & P3dx84);
	assign Q0dx84 = (W3dx84 | D4dx84);
	assign Lucx84 = (K4dx84 & R4dx84);
	assign R4dx84 = (Y4dx84 | F5dx84);
	assign K4dx84 = (M5dx84 & T5dx84);
	assign T5dx84 = (~(A6dx84 & H6dx84));
	assign A6dx84 = (~(O6dx84 & V6dx84));
	assign V6dx84 = (C7dx84 & J7dx84);
	assign J7dx84 = (~(Q7dx84 & X7dx84));
	assign Q7dx84 = (E8dx84 & L8dx84);
	assign L8dx84 = (~(S8dx84 & Z8dx84));
	assign S8dx84 = (Eobx84 ? G9dx84 : Q66w84);
	assign C7dx84 = (N9dx84 & U9dx84);
	assign N9dx84 = (~(Badx84 & Yrbx84));
	assign Badx84 = (~(W3dx84 | Hu2x84));
	assign O6dx84 = (Iadx84 & Padx84);
	assign Padx84 = (~(Wadx84 & Dbdx84));
	assign Dbdx84 = (Kbdx84 | Rbdx84);
	assign Rbdx84 = (~(Ybdx84 | Fcdx84));
	assign Kbdx84 = (Addx84 ? Tcdx84 : Mcdx84);
	assign Addx84 = (!Hddx84);
	assign Tcdx84 = (~(Eobx84 | Ba6w84));
	assign Iadx84 = (~(Oddx84 & Vddx84));
	assign Vddx84 = (~(Cedx84 & Jedx84));
	assign Jedx84 = (Qedx84 & Xedx84);
	assign Xedx84 = (Efdx84 | Lfdx84);
	assign Qedx84 = (~(Sfdx84 | Zfdx84));
	assign Sfdx84 = (Ggdx84 & Q66w84);
	assign Cedx84 = (Ngdx84 & Ugdx84);
	assign Ugdx84 = (Bhdx84 | Ihdx84);
	assign Ngdx84 = (~(Gwbx84 & Eobx84));
	assign M5dx84 = (~(Phdx84 & Whdx84));
	assign Whdx84 = (~(Didx84 & Kidx84));
	assign Kidx84 = (Ridx84 & Yidx84);
	assign Yidx84 = (~(Yrbx84 & Fjdx84));
	assign Fjdx84 = (~(Mjdx84 & Tjdx84));
	assign Tjdx84 = (Akdx84 | Hkdx84);
	assign Mjdx84 = (Okdx84 & Vkdx84);
	assign Okdx84 = (Cldx84 | D53x84);
	assign Ridx84 = (Jldx84 & Qldx84);
	assign Jldx84 = (~(Xldx84 & Emdx84));
	assign Emdx84 = (Hu2x84 & Lmdx84);
	assign Xldx84 = (Aq4w84 & Y6bx84);
	assign Didx84 = (Smdx84 & Zmdx84);
	assign Zmdx84 = (Gndx84 | Yybx84);
	assign Smdx84 = (~(Nndx84 & Undx84));
	assign Kq8x84 = (Bodx84 ? X473a4[23] : HWDATA[23]);
	assign Eq8x84 = (~(Iodx84 & Podx84));
	assign Podx84 = (Wodx84 & Dpdx84);
	assign Dpdx84 = (~(Kpdx84 & Qp63a4[31]));
	assign Wodx84 = (Rpdx84 & Ypdx84);
	assign Rpdx84 = (~(Fqdx84 & Mqdx84));
	assign Iodx84 = (Tqdx84 & Ardx84);
	assign Ardx84 = (~(Cr63a4[30] & Hrdx84));
	assign Tqdx84 = (~(Tk63a4[30] & Ordx84));
	assign Yp8x84 = (Csdx84 ? Km63a4[0] : Vrdx84);
	assign Vrdx84 = (~(Jsdx84 & Qsdx84));
	assign Qsdx84 = (Xsdx84 & Etdx84);
	assign Etdx84 = (~(Mw5w84 & Ltdx84));
	assign Xsdx84 = (~(Kr5w84 & Stdx84));
	assign Jsdx84 = (Ztdx84 & Gudx84);
	assign Gudx84 = (~(Y46w84 & Nudx84));
	assign Sp8x84 = (Bvdx84 ? Uudx84 : Eo5w84);
	assign Uudx84 = (~(Ivdx84 & Pvdx84));
	assign Pvdx84 = (~(Wvdx84 & Dwdx84));
	assign Ivdx84 = (Kwdx84 & Rwdx84);
	assign Rwdx84 = (~(Ywdx84 & Fxdx84));
	assign Kwdx84 = (Mxdx84 | Txdx84);
	assign Mp8x84 = (~(Aydx84 & Hydx84));
	assign Hydx84 = (Oydx84 & Vydx84);
	assign Vydx84 = (~(Czdx84 & Eo5w84));
	assign Oydx84 = (~(Jzdx84 & HADDR[30]));
	assign Aydx84 = (Qzdx84 & Xzdx84);
	assign Xzdx84 = (~(E0ex84 & Tk63a4[29]));
	assign Qzdx84 = (~(Cgaw84 & L0ex84));
	assign Gp8x84 = (Z0ex84 ? S0ex84 : P25w84);
	assign Z0ex84 = (HREADY & G1ex84);
	assign G1ex84 = (~(Mxdx84 & N1ex84));
	assign N1ex84 = (~(U1ex84 & B2ex84));
	assign B2ex84 = (Nndx84 | I2ex84);
	assign I2ex84 = (Vx2x84 & Bw2x84);
	assign U1ex84 = (P2ex84 & W2ex84);
	assign P2ex84 = (Kpdx84 | Fqdx84);
	assign S0ex84 = (~(D3ex84 & K3ex84));
	assign K3ex84 = (~(Qp63a4[0] & R3ex84));
	assign D3ex84 = (Y3ex84 & F4ex84);
	assign F4ex84 = (Mxdx84 | M4ex84);
	assign Y3ex84 = (T4ex84 | A5ex84);
	assign Ap8x84 = (~(H5ex84 & O5ex84));
	assign O5ex84 = (V5ex84 & C6ex84);
	assign C6ex84 = (~(J6ex84 & HRDATA[31]));
	assign V5ex84 = (Q6ex84 & X6ex84);
	assign X6ex84 = (~(G72x84 & E7ex84));
	assign Q6ex84 = (~(L7ex84 & HRDATA[15]));
	assign H5ex84 = (S7ex84 & Z7ex84);
	assign Z7ex84 = (~(Gc1x84 & G8ex84));
	assign S7ex84 = (J8cx84 | N8ex84);
	assign Uo8x84 = (~(U8ex84 & B9ex84));
	assign B9ex84 = (~(I9ex84 & HREADY));
	assign I9ex84 = (P9ex84 & W9ex84);
	assign P9ex84 = (~(Daex84 & Kaex84));
	assign Kaex84 = (Raex84 | Vx2x84);
	assign Daex84 = (Yaex84 & Hscx84);
	assign Yaex84 = (~(Fbex84 & Mbex84));
	assign U8ex84 = (Tbex84 | Acex84);
	assign Oo8x84 = (~(Hcex84 & Ocex84));
	assign Ocex84 = (Vcex84 & Cdex84);
	assign Cdex84 = (~(HRDATA[29] & J6ex84));
	assign Vcex84 = (Jdex84 & Qdex84);
	assign Qdex84 = (~(O32x84 & E7ex84));
	assign Jdex84 = (~(HRDATA[13] & L7ex84));
	assign Hcex84 = (Xdex84 & Eeex84);
	assign Eeex84 = (~(O81x84 & G8ex84));
	assign Xdex84 = (Leex84 | N8ex84);
	assign Io8x84 = (~(Seex84 & Zeex84));
	assign Zeex84 = (Gfex84 & Nfex84);
	assign Nfex84 = (~(Cr63a4[7] & Hrdx84));
	assign Gfex84 = (Ufex84 & Bgex84);
	assign Bgex84 = (Igex84 | Pgex84);
	assign Ufex84 = (~(Kpdx84 & Qp63a4[8]));
	assign Seex84 = (Wgex84 & Dhex84);
	assign Dhex84 = (~(Tk63a4[7] & Ordx84));
	assign Co8x84 = (~(Khex84 & Rhex84));
	assign Rhex84 = (Yhex84 & Fiex84);
	assign Fiex84 = (~(Kpdx84 & Qp63a4[30]));
	assign Yhex84 = (Miex84 & Ypdx84);
	assign Miex84 = (Igex84 | Txdx84);
	assign Khex84 = (Tiex84 & Ajex84);
	assign Ajex84 = (~(Cr63a4[29] & Hrdx84));
	assign Tiex84 = (~(Tk63a4[29] & Ordx84));
	assign Wn8x84 = (~(Hjex84 & Ojex84));
	assign Ojex84 = (Vjex84 | HREADY);
	assign Hjex84 = (Ckex84 & Jkex84);
	assign Ckex84 = (~(Qkex84 & Xkex84));
	assign Qn8x84 = (Elex84 & Llex84);
	assign Llex84 = (~(Slex84 | Zlex84));
	assign Elex84 = (IRQ[0] & Gmex84);
	assign Gmex84 = (~(Nmex84 & Umex84));
	assign Kn8x84 = (Aq4w84 ? Inex84 : Bnex84);
	assign Inex84 = (~(Pnex84 & Wnex84));
	assign Bnex84 = (~(Doex84 & Koex84));
	assign Koex84 = (Roex84 & Yoex84);
	assign Roex84 = (~(RXEV | TXEV));
	assign Doex84 = (Fpex84 & Mpex84);
	assign Fpex84 = (~(R83x84 & Tpex84));
	assign Tpex84 = (~(Aqex84 & Hqex84));
	assign Hqex84 = (Oqex84 & Vqex84);
	assign Vqex84 = (Crex84 & Jrex84);
	assign Jrex84 = (Qrex84 | Js3x84);
	assign Crex84 = (Xrex84 & Esex84);
	assign Esex84 = (~(Lsex84 & Ssex84));
	assign Lsex84 = (~(Zsex84 | Kf3x84));
	assign Xrex84 = (~(Gtex84 & Ntex84));
	assign Gtex84 = (HWDATA[28] & Utex84);
	assign Utex84 = (!Td3x84);
	assign Oqex84 = (Buex84 & Iuex84);
	assign Iuex84 = (Puex84 | Cc3x84);
	assign Buex84 = (~(Wuex84 & Dvex84));
	assign Dvex84 = (~(Kvex84 & Rvex84));
	assign Rvex84 = (Yvex84 & Fwex84);
	assign Fwex84 = (Mwex84 & Twex84);
	assign Twex84 = (Axex84 & Hxex84);
	assign Hxex84 = (~(HWDATA[6] | HWDATA[7]));
	assign Axex84 = (~(HWDATA[4] | HWDATA[5]));
	assign Mwex84 = (~(Oxex84 | HWDATA[28]));
	assign Oxex84 = (HWDATA[29] | HWDATA[30]);
	assign Yvex84 = (Vxex84 & Cyex84);
	assign Cyex84 = (Jyex84 & Qyex84);
	assign Qyex84 = (~(HWDATA[26] | HWDATA[27]));
	assign Jyex84 = (~(HWDATA[24] | HWDATA[25]));
	assign Vxex84 = (Xyex84 & Ezex84);
	assign Xyex84 = (~(Lzex84 | Szex84));
	assign Kvex84 = (Zzex84 & G0fx84);
	assign G0fx84 = (N0fx84 & U0fx84);
	assign U0fx84 = (B1fx84 & I1fx84);
	assign I1fx84 = (~(HWDATA[11] | HWDATA[10]));
	assign B1fx84 = (~(HWDATA[13] | HWDATA[12]));
	assign N0fx84 = (P1fx84 & W1fx84);
	assign P1fx84 = (~(HWDATA[15] | HWDATA[14]));
	assign Zzex84 = (D2fx84 & K2fx84);
	assign K2fx84 = (R2fx84 & Y2fx84);
	assign Y2fx84 = (~(HWDATA[18] | HWDATA[17]));
	assign R2fx84 = (~(HWDATA[20] | HWDATA[19]));
	assign D2fx84 = (F3fx84 & M3fx84);
	assign F3fx84 = (~(HWDATA[8] | HWDATA[21]));
	assign Aqex84 = (T3fx84 & A4fx84);
	assign A4fx84 = (H4fx84 & O4fx84);
	assign O4fx84 = (~(Ye63a4 & V4fx84));
	assign V4fx84 = (!K873a4[1]);
	assign Ye63a4 = (~(C5fx84 & J5fx84));
	assign J5fx84 = (~(IRQ[1] & Q5fx84));
	assign C5fx84 = (~(X5fx84 & E6fx84));
	assign X5fx84 = (L6fx84 & S6fx84);
	assign S6fx84 = (Z6fx84 | K873a4[1]);
	assign L6fx84 = (G7fx84 | N7fx84);
	assign H4fx84 = (U7fx84 & B8fx84);
	assign B8fx84 = (~(Mf63a4 & I8fx84));
	assign I8fx84 = (!K873a4[3]);
	assign Mf63a4 = (~(P8fx84 & W8fx84));
	assign W8fx84 = (~(IRQ[3] & D9fx84));
	assign P8fx84 = (~(K9fx84 & R9fx84));
	assign R9fx84 = (Y9fx84 | Yoex84);
	assign K9fx84 = (Fafx84 & Mafx84);
	assign Mafx84 = (Tafx84 | K873a4[3]);
	assign Fafx84 = (Abfx84 | N7fx84);
	assign U7fx84 = (~(Ff63a4 & Hbfx84));
	assign Hbfx84 = (!K873a4[0]);
	assign Ff63a4 = (~(Obfx84 & Vbfx84));
	assign Vbfx84 = (~(IRQ[0] & Slex84));
	assign Slex84 = (X54x84 & Ccfx84);
	assign Obfx84 = (~(Jcfx84 & Ccfx84));
	assign Ccfx84 = (~(Umex84 & Qcfx84));
	assign Jcfx84 = (Xcfx84 & Edfx84);
	assign Edfx84 = (Zlex84 | K873a4[0]);
	assign Zlex84 = (HWDATA[0] & Wuex84);
	assign Xcfx84 = (Ldfx84 | N7fx84);
	assign T3fx84 = (Sdfx84 & Zdfx84);
	assign Zdfx84 = (Gefx84 | K873a4[2]);
	assign Gefx84 = (!Re63a4);
	assign Re63a4 = (Nefx84 & Uefx84);
	assign Uefx84 = (~(Bffx84 & Iffx84));
	assign Iffx84 = (~(IRQ[2] & Pffx84));
	assign Bffx84 = (Wffx84 & Dgfx84);
	assign Wffx84 = (~(K873a4[2] & Kgfx84));
	assign Kgfx84 = (N7fx84 | Rgfx84);
	assign N7fx84 = (~(Ygfx84 & Fhfx84));
	assign Sdfx84 = (~(Yi3x84 & Mhfx84));
	assign Yi3x84 = (Thfx84 & Aifx84);
	assign Aifx84 = (~(Hifx84 & Oifx84));
	assign Oifx84 = (~(NMI & Vifx84));
	assign Hifx84 = (Cjfx84 & Mhfx84);
	assign En8x84 = (~(Jjfx84 & Qjfx84));
	assign Qjfx84 = (Xjfx84 & Ekfx84);
	assign Ekfx84 = (~(Czdx84 & Up5w84));
	assign Xjfx84 = (~(Jzdx84 & HADDR[31]));
	assign Jjfx84 = (Lkfx84 & Skfx84);
	assign Skfx84 = (~(E0ex84 & Tk63a4[30]));
	assign Lkfx84 = (~(Yhaw84 & L0ex84));
	assign Ym8x84 = (Zkfx84 | Glfx84);
	assign Zkfx84 = (Ulfx84 ? Nlfx84 : Ce1x84);
	assign Sm8x84 = (Bmfx84 | Imfx84);
	assign Imfx84 = (N8ex84 ? Pmfx84 : W05w84);
	assign Pmfx84 = (~(Wmfx84 | Dnfx84));
	assign Bmfx84 = (~(Knfx84 & Rnfx84));
	assign Rnfx84 = (~(C92x84 & E7ex84));
	assign Knfx84 = (~(Ce1x84 & G8ex84));
	assign Mm8x84 = (Ynfx84 & Fofx84);
	assign Fofx84 = (~(Mofx84 & Tofx84));
	assign Tofx84 = (Apfx84 & Hpfx84);
	assign Apfx84 = (~(Opfx84 & Vpfx84));
	assign Vpfx84 = (~(Cqfx84 & Jqfx84));
	assign Jqfx84 = (Qqfx84 & Xqfx84);
	assign Qqfx84 = (Erfx84 & Lrfx84);
	assign Cqfx84 = (Srfx84 & Zrfx84);
	assign Srfx84 = (~(Fn2x84 & Gsfx84));
	assign Gsfx84 = (~(Mw5w84 & Nsfx84));
	assign Nsfx84 = (Kr5w84 | Ct5w84);
	assign Opfx84 = (Yk5w84 | Usfx84);
	assign Usfx84 = (Yybx84 & V55w84);
	assign Mofx84 = (Btfx84 & HREADY);
	assign Btfx84 = (Kr5w84 ? Ptfx84 : Itfx84);
	assign Ptfx84 = (Wtfx84 | Qtcx84);
	assign Itfx84 = (~(Dufx84 & Kufx84));
	assign Kufx84 = (~(Ambx84 | D4dx84));
	assign Dufx84 = (~(Rufx84 | Yufx84));
	assign Ynfx84 = (~(Fvfx84 & Mvfx84));
	assign Mvfx84 = (~(HREADY & Hpfx84));
	assign Hpfx84 = (~(Tvfx84 & Awfx84));
	assign Awfx84 = (Hwfx84 & Owfx84);
	assign Owfx84 = (~(Vwfx84 | Cxfx84));
	assign Hwfx84 = (Jxfx84 & Qxfx84);
	assign Tvfx84 = (Xxfx84 & Eyfx84);
	assign Eyfx84 = (Lyfx84 & Syfx84);
	assign Syfx84 = (~(Zyfx84 & Pxbx84));
	assign Zyfx84 = (~(Gzfx84 | Vx2x84));
	assign Lyfx84 = (~(Nzfx84 & Uzfx84));
	assign Uzfx84 = (~(B0gx84 & I0gx84));
	assign I0gx84 = (~(P0gx84 & Gpbx84));
	assign Xxfx84 = (W0gx84 & D1gx84);
	assign W0gx84 = (Tq2x84 ? R1gx84 : K1gx84);
	assign R1gx84 = (~(Y1gx84 & Zo2x84));
	assign K1gx84 = (~(F2gx84 & M2gx84));
	assign M2gx84 = (~(Lrfx84 & T2gx84));
	assign T2gx84 = (Gzfx84 | Gz4w84);
	assign Gm8x84 = (~(A3gx84 & H3gx84));
	assign H3gx84 = (O3gx84 & V3gx84);
	assign V3gx84 = (~(Czdx84 & Hj5w84));
	assign O3gx84 = (~(Jzdx84 & HADDR[9]));
	assign A3gx84 = (C4gx84 & J4gx84);
	assign J4gx84 = (~(Tk63a4[8] & E0ex84));
	assign C4gx84 = (~(Jd9w84 & L0ex84));
	assign Am8x84 = (X4gx84 ? U9xw84 : Q4gx84);
	assign Ul8x84 = (X4gx84 ? Qbxw84 : E5gx84);
	assign Ol8x84 = (X4gx84 ? Psvw84 : L5gx84);
	assign Il8x84 = (Z5gx84 ? S5gx84 : Yk5w84);
	assign Z5gx84 = (HREADY & G6gx84);
	assign G6gx84 = (~(N6gx84 & U6gx84));
	assign U6gx84 = (~(B7gx84 & I7gx84));
	assign I7gx84 = (Wl6w84 & P7gx84);
	assign B7gx84 = (~(W7gx84 | D8gx84));
	assign N6gx84 = (~(Yybx84 | Qcfx84));
	assign S5gx84 = (~(K8gx84 & R8gx84));
	assign R8gx84 = (~(P7gx84 & Y8gx84));
	assign K8gx84 = (~(Bg5w84 & V55w84));
	assign Cl8x84 = (X4gx84 ? Kuvw84 : F9gx84);
	assign Wk8x84 = (~(M9gx84 & T9gx84));
	assign T9gx84 = (Aagx84 & Hagx84);
	assign Hagx84 = (~(Cr63a4[22] & Hrdx84));
	assign Aagx84 = (Oagx84 & Vagx84);
	assign Vagx84 = (Igex84 | Cbgx84);
	assign Oagx84 = (~(Qp63a4[23] & Kpdx84));
	assign M9gx84 = (Jbgx84 & Qbgx84);
	assign Qbgx84 = (~(Tk63a4[22] & Ordx84));
	assign Qk8x84 = (X4gx84 ? Wwww84 : Xbgx84);
	assign Kk8x84 = (~(Ecgx84 & Lcgx84));
	assign Lcgx84 = (Scgx84 | HREADY);
	assign Ecgx84 = (Zcgx84 & Jkex84);
	assign Zcgx84 = (~(Qkex84 & Gdgx84));
	assign Gdgx84 = (HADDR[2] | HADDR[7]);
	assign Ek8x84 = (~(Ndgx84 & Udgx84));
	assign Udgx84 = (~(T14x84 & Wpcx84));
	assign Ndgx84 = (Begx84 & Jkex84);
	assign Begx84 = (~(Qkex84 & Iegx84));
	assign Iegx84 = (HADDR[3] | HADDR[5]);
	assign Yj8x84 = (~(Pegx84 & Wegx84));
	assign Wegx84 = (Dfgx84 | HREADY);
	assign Pegx84 = (Kfgx84 & Jkex84);
	assign Kfgx84 = (~(Qkex84 & Rfgx84));
	assign Rfgx84 = (~(HADDR[10] ^ Yfgx84));
	assign Sj8x84 = (~(Fggx84 & Mggx84));
	assign Mggx84 = (~(Zx3x84 & Wpcx84));
	assign Fggx84 = (Tggx84 & Jkex84);
	assign Jkex84 = (~(Qkex84 & Ahgx84));
	assign Ahgx84 = (~(Hhgx84 & Ohgx84));
	assign Ohgx84 = (Vhgx84 & Cigx84);
	assign Cigx84 = (Jigx84 & Qigx84);
	assign Qigx84 = (~(Xigx84 | HADDR[26]));
	assign Xigx84 = (HADDR[27] | HADDR[6]);
	assign Jigx84 = (~(HADDR[24] | HADDR[25]));
	assign Vhgx84 = (Ejgx84 & Ljgx84);
	assign Ljgx84 = (~(Sjgx84 | HADDR[21]));
	assign Sjgx84 = (HADDR[22] | HADDR[23]);
	assign Ejgx84 = (~(HADDR[19] | HADDR[20]));
	assign Hhgx84 = (Zjgx84 & Gkgx84);
	assign Gkgx84 = (Nkgx84 & Ukgx84);
	assign Ukgx84 = (~(Blgx84 | HADDR[16]));
	assign Blgx84 = (HADDR[17] | HADDR[18]);
	assign Nkgx84 = (HSIZE[1] & Ilgx84);
	assign Ilgx84 = (!HADDR[12]);
	assign Zjgx84 = (Plgx84 & Wlgx84);
	assign Wlgx84 = (HADDR[14] & HADDR[15]);
	assign Plgx84 = (Dmgx84 & HADDR[13]);
	assign Dmgx84 = (~(Kmgx84 & Rmgx84));
	assign Rmgx84 = (~(Ymgx84 & Fngx84));
	assign Fngx84 = (Mngx84 & Tngx84);
	assign Tngx84 = (!HADDR[5]);
	assign Mngx84 = (~(HADDR[7] | HADDR[9]));
	assign Ymgx84 = (Aogx84 & Hogx84);
	assign Hogx84 = (~(Oogx84 & Vogx84));
	assign Oogx84 = (~(HADDR[10] | HADDR[4]));
	assign Aogx84 = (HADDR[11] ? Cpgx84 : Xkex84);
	assign Cpgx84 = (Jpgx84 & Vogx84);
	assign Vogx84 = (Yfgx84 | HADDR[2]);
	assign Yfgx84 = (!HADDR[3]);
	assign Jpgx84 = (~(Qpgx84 | Xkex84));
	assign Kmgx84 = (~(Xpgx84 & Eqgx84));
	assign Eqgx84 = (Lqgx84 & Sqgx84);
	assign Sqgx84 = (!HADDR[2]);
	assign Lqgx84 = (~(HADDR[3] | HADDR[4]));
	assign Xpgx84 = (Zqgx84 & Grgx84);
	assign Grgx84 = (HADDR[8] ^ HADDR[9]);
	assign Zqgx84 = (Qpgx84 ? Urgx84 : Nrgx84);
	assign Qpgx84 = (!HADDR[10]);
	assign Urgx84 = (~(HADDR[11] | HADDR[5]));
	assign Nrgx84 = (Bsgx84 & HADDR[11]);
	assign Bsgx84 = (~(Xkex84 | HADDR[7]));
	assign Xkex84 = (!HADDR[8]);
	assign Tggx84 = (Isgx84 | HADDR[4]);
	assign Isgx84 = (!Qkex84);
	assign Mj8x84 = (~(Psgx84 & Wsgx84));
	assign Wsgx84 = (~(R673a4[0] & Dtgx84));
	assign Dtgx84 = (Ldfx84 | Ktgx84);
	assign Psgx84 = (Rtgx84 | Ldfx84);
	assign Ldfx84 = (!HWDATA[0]);
	assign Gj8x84 = (~(Ytgx84 & Fugx84));
	assign Fugx84 = (~(Dj0x84 & Yoex84));
	assign Aj8x84 = (~(Mugx84 & Tugx84));
	assign Tugx84 = (Avgx84 | Hvgx84);
	assign Hvgx84 = (C45w84 ? Vvgx84 : Ovgx84);
	assign Ovgx84 = (Hscx84 | Cwgx84);
	assign Avgx84 = (Jwgx84 | H6dx84);
	assign Mugx84 = (~(Nx4w84 & Qwgx84));
	assign Ui8x84 = (~(Xwgx84 & Exgx84));
	assign Exgx84 = (Lxgx84 & Sxgx84);
	assign Sxgx84 = (~(Kpdx84 & Qp63a4[1]));
	assign Lxgx84 = (Zxgx84 & Ypdx84);
	assign Zxgx84 = (Igex84 | Gygx84);
	assign Xwgx84 = (Nygx84 & Uygx84);
	assign Uygx84 = (~(Cr63a4[0] & Hrdx84));
	assign Nygx84 = (Bzgx84 | Izgx84);
	assign Oi8x84 = (Qkex84 ? HWRITE : Pzgx84);
	assign Qkex84 = (Wzgx84 & D0hx84);
	assign D0hx84 = (K0hx84 & R0hx84);
	assign R0hx84 = (~(Y0hx84 | HADDR[28]));
	assign K0hx84 = (~(F1hx84 | M1hx84));
	assign Wzgx84 = (~(T1hx84 | A2hx84));
	assign T1hx84 = (~(H2hx84 & O2hx84));
	assign Pzgx84 = (V2hx84 & C3hx84);
	assign Ii8x84 = (~(J3hx84 & Q3hx84));
	assign Q3hx84 = (~(R673a4[3] & X3hx84));
	assign X3hx84 = (Abfx84 | Ktgx84);
	assign J3hx84 = (Rtgx84 | Abfx84);
	assign Abfx84 = (!HWDATA[3]);
	assign Ci8x84 = (~(E4hx84 & L4hx84));
	assign L4hx84 = (~(R673a4[2] & S4hx84));
	assign S4hx84 = (Rgfx84 | Ktgx84);
	assign E4hx84 = (Rtgx84 | Rgfx84);
	assign Rgfx84 = (!HWDATA[2]);
	assign Wh8x84 = (~(Z4hx84 & G5hx84));
	assign G5hx84 = (~(R673a4[1] & N5hx84));
	assign N5hx84 = (G7fx84 | Ktgx84);
	assign Ktgx84 = (Rtgx84 & U5hx84);
	assign U5hx84 = (~(B6hx84 & Fhfx84));
	assign B6hx84 = (In4w84 & I6hx84);
	assign Z4hx84 = (Rtgx84 | G7fx84);
	assign G7fx84 = (!HWDATA[1]);
	assign Rtgx84 = (~(C3hx84 & I6hx84));
	assign Qh8x84 = (P6hx84 ? Qm3x84 : HWDATA[2]);
	assign Kh8x84 = (P6hx84 ? Oo3x84 : HWDATA[1]);
	assign Eh8x84 = (P6hx84 ? Mq3x84 : HWDATA[0]);
	assign P6hx84 = (~(W6hx84 & In4w84));
	assign Yg8x84 = (Bodx84 ? X473a4[22] : Lzex84);
	assign Sg8x84 = (Bodx84 ? X473a4[21] : HWDATA[21]);
	assign Mg8x84 = (Bodx84 ? X473a4[20] : HWDATA[20]);
	assign Gg8x84 = (Bodx84 ? X473a4[19] : HWDATA[19]);
	assign Ag8x84 = (Bodx84 ? X473a4[18] : HWDATA[18]);
	assign Uf8x84 = (Bodx84 ? X473a4[17] : HWDATA[17]);
	assign Of8x84 = (Bodx84 ? X473a4[16] : HWDATA[16]);
	assign If8x84 = (Bodx84 ? X473a4[15] : HWDATA[15]);
	assign Cf8x84 = (Bodx84 ? X473a4[14] : HWDATA[14]);
	assign We8x84 = (Bodx84 ? X473a4[13] : HWDATA[13]);
	assign Qe8x84 = (Bodx84 ? X473a4[12] : HWDATA[12]);
	assign Ke8x84 = (Bodx84 ? X473a4[11] : HWDATA[11]);
	assign Ee8x84 = (Bodx84 ? X473a4[10] : HWDATA[10]);
	assign Yd8x84 = (Bodx84 ? X473a4[9] : HWDATA[9]);
	assign Sd8x84 = (Bodx84 ? X473a4[8] : HWDATA[8]);
	assign Md8x84 = (Bodx84 ? X473a4[7] : HWDATA[7]);
	assign Gd8x84 = (Bodx84 ? X473a4[6] : HWDATA[6]);
	assign Ad8x84 = (Bodx84 ? X473a4[5] : HWDATA[5]);
	assign Uc8x84 = (Bodx84 ? X473a4[4] : HWDATA[4]);
	assign Bodx84 = (!D7hx84);
	assign Oc8x84 = (D7hx84 ? HWDATA[3] : X473a4[3]);
	assign Ic8x84 = (D7hx84 ? HWDATA[2] : X473a4[2]);
	assign Cc8x84 = (D7hx84 ? HWDATA[1] : X473a4[1]);
	assign Wb8x84 = (D7hx84 ? HWDATA[0] : X473a4[0]);
	assign D7hx84 = (K7hx84 & R7hx84);
	assign K7hx84 = (Fhfx84 & In4w84);
	assign Qb8x84 = (Y7hx84 ? Nz63a4[0] : HWDATA[6]);
	assign Kb8x84 = (Y7hx84 ? Nz63a4[1] : HWDATA[7]);
	assign Eb8x84 = (Y7hx84 ? Nz63a4[2] : HWDATA[14]);
	assign Ya8x84 = (Y7hx84 ? Nz63a4[3] : HWDATA[15]);
	assign Y7hx84 = (!F8hx84);
	assign Sa8x84 = (F8hx84 ? Lzex84 : Nz63a4[4]);
	assign Ma8x84 = (F8hx84 ? HWDATA[23] : Nz63a4[5]);
	assign Ga8x84 = (F8hx84 ? HWDATA[30] : Nz63a4[6]);
	assign Aa8x84 = (F8hx84 ? Szex84 : Nz63a4[7]);
	assign F8hx84 = (Ygfx84 & M8hx84);
	assign Ygfx84 = (T8hx84 & In4w84);
	assign U98x84 = (A9hx84 ? HWDATA[1] : Lo4w84);
	assign O98x84 = (A9hx84 ? HWDATA[2] : Y63x84);
	assign A9hx84 = (!H9hx84);
	assign I98x84 = (H9hx84 ? R83x84 : HWDATA[4]);
	assign H9hx84 = (~(O9hx84 & M8hx84));
	assign O9hx84 = (V2hx84 & In4w84);
	assign C98x84 = (V9hx84 ? Szex84 : Xx63a4[1]);
	assign W88x84 = (V9hx84 ? HWDATA[30] : Xx63a4[0]);
	assign V9hx84 = (Cahx84 & In4w84);
	assign Q88x84 = (Jahx84 ? Hw63a4[1] : HWDATA[23]);
	assign K88x84 = (Jahx84 ? Hw63a4[0] : Lzex84);
	assign E88x84 = (Jahx84 ? D373a4[1] : Szex84);
	assign Y78x84 = (Jahx84 ? D373a4[0] : HWDATA[30]);
	assign Jahx84 = (~(Qahx84 & Xahx84));
	assign Xahx84 = (Ebhx84 & I6hx84);
	assign Qahx84 = (T14x84 & In4w84);
	assign S78x84 = (~(Lbhx84 & Sbhx84));
	assign Sbhx84 = (~(Zbhx84 & Vk3x84));
	assign Zbhx84 = (~(Gchx84 | Nchx84));
	assign Gchx84 = (~(Uchx84 | In4w84));
	assign Uchx84 = (!W6hx84);
	assign Lbhx84 = (~(Bdhx84 & Idhx84));
	assign Bdhx84 = (Pdhx84 & Pu63a4[0]);
	assign M78x84 = (X4gx84 ? Uqvw84 : Wdhx84);
	assign G78x84 = (Dehx84 | Kehx84);
	assign Dehx84 = (HREADY ? Rehx84 : Nr4w84);
	assign Rehx84 = (~(Yehx84 | Ffhx84));
	assign Yehx84 = (Mfhx84 & Tfhx84);
	assign Tfhx84 = (~(Aghx84 & Hghx84));
	assign Aghx84 = (~(Wbcx84 | Oghx84));
	assign Mfhx84 = (~(P7gx84 & Vghx84));
	assign A78x84 = (~(Chhx84 & Jhhx84));
	assign Jhhx84 = (Qhhx84 & Xhhx84);
	assign Xhhx84 = (~(Kpdx84 & Qp63a4[29]));
	assign Qhhx84 = (Eihx84 & Ypdx84);
	assign Eihx84 = (Igex84 | Lihx84);
	assign Chhx84 = (Sihx84 & Zihx84);
	assign Zihx84 = (~(Cr63a4[28] & Hrdx84));
	assign Sihx84 = (~(Tk63a4[28] & Ordx84));
	assign U68x84 = (Gjhx84 ? Khsw84 : Wdhx84);
	assign O68x84 = (Gjhx84 ? Fjsw84 : L5gx84);
	assign I68x84 = (Gjhx84 ? Alsw84 : F9gx84);
	assign C68x84 = (Gjhx84 ? Busw84 : Njhx84);
	assign W58x84 = (~(Ujhx84 & Bkhx84));
	assign Bkhx84 = (~(Ntex84 & HWDATA[28]));
	assign Ujhx84 = (~(Ikhx84 & Td3x84));
	assign Ikhx84 = (Pkhx84 & Wkhx84);
	assign Wkhx84 = (~(Ntex84 & HWDATA[27]));
	assign Pkhx84 = (~(Dlhx84 & Qcfx84));
	assign Q58x84 = (~(Klhx84 & Rlhx84));
	assign Rlhx84 = (Ylhx84 & Fmhx84);
	assign Fmhx84 = (~(Qp63a4[3] & Kpdx84));
	assign Ylhx84 = (Mmhx84 & Ypdx84);
	assign Mmhx84 = (Igex84 | Tmhx84);
	assign Klhx84 = (Anhx84 & Hnhx84);
	assign Hnhx84 = (~(Cr63a4[2] & Hrdx84));
	assign Anhx84 = (~(Tk63a4[2] & Ordx84));
	assign K58x84 = (~(Onhx84 & Vnhx84));
	assign Vnhx84 = (Cohx84 & Johx84);
	assign Johx84 = (~(J6ex84 & HRDATA[16]));
	assign Cohx84 = (Qohx84 & Xohx84);
	assign Xohx84 = (~(Yf1x84 & E7ex84));
	assign Qohx84 = (~(L7ex84 & HRDATA[0]));
	assign Onhx84 = (Ephx84 & Lphx84);
	assign Lphx84 = (~(Yk0x84 & G8ex84));
	assign Ephx84 = (Sphx84 | N8ex84);
	assign E58x84 = (Gqhx84 ? Zphx84 : Si6w84);
	assign Zphx84 = (~(Nqhx84 & Uqhx84));
	assign Uqhx84 = (Brhx84 & Irhx84);
	assign Irhx84 = (Prhx84 & Wrhx84);
	assign Wrhx84 = (~(Phdx84 & Dshx84));
	assign Dshx84 = (~(Kshx84 & Rshx84));
	assign Rshx84 = (Yshx84 | Fthx84);
	assign Prhx84 = (Mthx84 & Tthx84);
	assign Tthx84 = (~(Auhx84 & Huhx84));
	assign Auhx84 = (~(Ouhx84 | Ba6w84));
	assign Mthx84 = (~(Vuhx84 & Cvhx84));
	assign Vuhx84 = (Jvhx84 ^ Qvhx84);
	assign Brhx84 = (Xvhx84 & Ewhx84);
	assign Ewhx84 = (~(Lwhx84 & Yk0x84));
	assign Xvhx84 = (~(O16w84 & Swhx84));
	assign Nqhx84 = (Zwhx84 & Gxhx84);
	assign Gxhx84 = (Nxhx84 & Uxhx84);
	assign Uxhx84 = (Sphx84 | Byhx84);
	assign Nxhx84 = (Iyhx84 | Si6w84);
	assign Zwhx84 = (~(Pyhx84 | Wyhx84));
	assign Wyhx84 = (!Dzhx84);
	assign Pyhx84 = (Hu2x84 ? Qvax84 : Kzhx84);
	assign Kzhx84 = (Rzhx84 & Yzhx84);
	assign Y48x84 = (Fdcx84 ? F0ix84 : Ap6w84);
	assign Fdcx84 = (HREADY & M0ix84);
	assign M0ix84 = (~(T0ix84 & A1ix84));
	assign A1ix84 = (H1ix84 & O1ix84);
	assign O1ix84 = (~(V1ix84 & C2ix84));
	assign H1ix84 = (J2ix84 & Q2ix84);
	assign Q2ix84 = (~(X2ix84 & E3ix84));
	assign X2ix84 = (Nacx84 & Pxbx84);
	assign J2ix84 = (~(L3ix84 & S3ix84));
	assign T0ix84 = (Z3ix84 & G4ix84);
	assign G4ix84 = (~(Iqbx84 & N4ix84));
	assign F0ix84 = (~(U4ix84 & B5ix84));
	assign B5ix84 = (I5ix84 & P5ix84);
	assign P5ix84 = (W5ix84 & D6ix84);
	assign D6ix84 = (~(K6ix84 & R6ix84));
	assign R6ix84 = (P3dx84 ^ Y6ix84);
	assign Y6ix84 = (I3dx84 & Ln6w84);
	assign P3dx84 = (~(D8gx84 | J13x84));
	assign K6ix84 = (F7ix84 & M7ix84);
	assign W5ix84 = (T7ix84 & A8ix84);
	assign I5ix84 = (H8ix84 & O8ix84);
	assign O8ix84 = (~(V8ix84 & Ap6w84));
	assign V8ix84 = (Lgcx84 & C9ix84);
	assign Lgcx84 = (~(J9ix84 & Q9ix84));
	assign Q9ix84 = (X9ix84 & Tlbx84);
	assign Tlbx84 = (~(Phdx84 & Eaix84));
	assign Eaix84 = (Zo2x84 | Laix84);
	assign X9ix84 = (Erfx84 & Saix84);
	assign J9ix84 = (Zaix84 & Gbix84);
	assign Gbix84 = (~(Nacx84 & Mlbx84));
	assign Zaix84 = (Nbix84 | Pqbx84);
	assign H8ix84 = (~(I86w84 & Ubix84));
	assign Ubix84 = (~(Bcix84 & Icix84));
	assign Icix84 = (~(Pcix84 & V1ix84));
	assign U4ix84 = (Wcix84 & Ddix84);
	assign Ddix84 = (Kdix84 & Rdix84);
	assign Rdix84 = (~(Es0x84 & Encx84));
	assign Encx84 = (Dj0x84 & Ydix84);
	assign Ydix84 = (~(Feix84 & Meix84));
	assign Feix84 = (~(Teix84 | Afix84));
	assign Kdix84 = (Hfix84 & Ofix84);
	assign Ofix84 = (Rufx84 | Qfcx84);
	assign Qfcx84 = (Mebx84 & Vfix84);
	assign Vfix84 = (Cgix84 | Ouhx84);
	assign Hfix84 = (~(Ey5w84 & Picx84));
	assign Picx84 = (~(Oecx84 & Cfcx84));
	assign Oecx84 = (Jgix84 & Qgix84);
	assign Qgix84 = (Xgix84 & Ehix84);
	assign Ehix84 = (~(Lhix84 & Shix84));
	assign Lhix84 = (~(Ouhx84 | Nd6w84));
	assign Jgix84 = (Zhix84 & Giix84);
	assign Giix84 = (Niix84 | Qtcx84);
	assign Wcix84 = (Uiix84 & Bjix84);
	assign Bjix84 = (Lncx84 | Wcbx84);
	assign S48x84 = (~(Ijix84 & Pjix84));
	assign Pjix84 = (~(Wjix84 & M1hx84));
	assign Wjix84 = (H2hx84 & Dkix84);
	assign Ijix84 = (~(Kkix84 & Wpcx84));
	assign Kkix84 = (~(H6dx84 & Rkix84));
	assign Rkix84 = (~(HRESP & Ykix84));
	assign Ykix84 = (~(Flix84 & Mlix84));
	assign Mlix84 = (Tlix84 & Amix84);
	assign Amix84 = (Hmix84 & Omix84);
	assign Omix84 = (~(Vmix84 & Cnix84));
	assign Cnix84 = (~(Jnix84 | Bw2x84));
	assign Vmix84 = (~(Fthx84 | Ambx84));
	assign Hmix84 = (Qnix84 & Nbix84);
	assign Tlix84 = (Xnix84 & Eoix84);
	assign Eoix84 = (~(Loix84 & Soix84));
	assign Loix84 = (~(N4ix84 | Tq2x84));
	assign Xnix84 = (~(Zoix84 & Gpix84));
	assign Flix84 = (Npix84 & Upix84);
	assign Upix84 = (Bqix84 & Iqix84);
	assign Iqix84 = (Pqix84 | Pqbx84);
	assign Bqix84 = (Wqix84 & Drix84);
	assign Drix84 = (~(Krix84 & Rrix84));
	assign Rrix84 = (~(Yrix84 & Fsix84));
	assign Fsix84 = (~(Msix84 & F2gx84));
	assign Msix84 = (~(Tsix84 | Hu2x84));
	assign Wqix84 = (~(Atix84 & Htix84));
	assign Htix84 = (~(Otix84 & Vtix84));
	assign Vtix84 = (Cuix84 | Tsix84);
	assign Otix84 = (Juix84 & Quix84);
	assign Juix84 = (~(Xuix84 & Drbx84));
	assign Xuix84 = (~(Evix84 | Fn2x84));
	assign Npix84 = (Lvix84 & Svix84);
	assign Svix84 = (~(Zvix84 & Gwix84));
	assign Lvix84 = (~(Nwix84 & Uwix84));
	assign M48x84 = (~(Bxix84 & Ixix84));
	assign Ixix84 = (Pxix84 & Wxix84);
	assign Wxix84 = (~(Qp63a4[7] & Kpdx84));
	assign Pxix84 = (Dyix84 & Ypdx84);
	assign Dyix84 = (~(Fqdx84 & Kyix84));
	assign Bxix84 = (Ryix84 & Yyix84);
	assign Yyix84 = (~(Cr63a4[6] & Hrdx84));
	assign Ryix84 = (~(Tk63a4[6] & Ordx84));
	assign G48x84 = (~(Fzix84 & Mzix84));
	assign Mzix84 = (Tzix84 & A0jx84);
	assign A0jx84 = (~(Cr63a4[14] & Hrdx84));
	assign Tzix84 = (H0jx84 & O0jx84);
	assign O0jx84 = (Igex84 | V0jx84);
	assign H0jx84 = (~(Qp63a4[15] & Kpdx84));
	assign Fzix84 = (Wgex84 & C1jx84);
	assign C1jx84 = (~(Tk63a4[14] & Ordx84));
	assign A48x84 = (J1jx84 | Glfx84);
	assign J1jx84 = (X1jx84 ? Gc1x84 : Q1jx84);
	assign Q1jx84 = (Dnfx84 & HRDATA[15]);
	assign Dnfx84 = (!Nlfx84);
	assign U38x84 = (~(E2jx84 & L2jx84));
	assign L2jx84 = (~(S2jx84 & HRDATA[14]));
	assign E2jx84 = (~(Ka1x84 & X1jx84));
	assign O38x84 = (~(Z2jx84 & G3jx84));
	assign G3jx84 = (~(S2jx84 & HRDATA[13]));
	assign Z2jx84 = (N3jx84 & Ytgx84);
	assign N3jx84 = (~(O81x84 & U3jx84));
	assign U3jx84 = (~(Ulfx84 & B4jx84));
	assign B4jx84 = (~(Dj0x84 & I4jx84));
	assign I4jx84 = (~(P4jx84 & W4jx84));
	assign W4jx84 = (!S61x84);
	assign I38x84 = (D5jx84 | K5jx84);
	assign K5jx84 = (S61x84 ? R5jx84 : P4jx84);
	assign R5jx84 = (~(Ulfx84 & Y5jx84));
	assign Y5jx84 = (P4jx84 | F6jx84);
	assign D5jx84 = (~(M6jx84 & Ytgx84));
	assign M6jx84 = (~(HRDATA[12] & S2jx84));
	assign C38x84 = (~(T6jx84 & A7jx84));
	assign A7jx84 = (~(P4jx84 | H7jx84));
	assign H7jx84 = (!Ytgx84);
	assign P4jx84 = (~(O7jx84 | W41x84));
	assign T6jx84 = (V7jx84 & C8jx84);
	assign C8jx84 = (~(W41x84 & J8jx84));
	assign J8jx84 = (~(Ulfx84 & Q8jx84));
	assign Q8jx84 = (~(O7jx84 & Glfx84));
	assign V7jx84 = (~(S2jx84 & HRDATA[11]));
	assign W28x84 = (~(X8jx84 & E9jx84));
	assign E9jx84 = (O7jx84 & Ytgx84);
	assign O7jx84 = (~(L9jx84 & S9jx84));
	assign L9jx84 = (~(A31x84 | F11x84));
	assign X8jx84 = (Z9jx84 & Gajx84);
	assign Gajx84 = (~(A31x84 & Najx84));
	assign Najx84 = (~(Uajx84 & Bbjx84));
	assign Bbjx84 = (~(F11x84 & Glfx84));
	assign Z9jx84 = (~(S2jx84 & HRDATA[10]));
	assign Q28x84 = (~(Ibjx84 & Pbjx84));
	assign Pbjx84 = (F11x84 ? Uajx84 : Wbjx84);
	assign Uajx84 = (Ulfx84 & Dcjx84);
	assign Dcjx84 = (S9jx84 | F6jx84);
	assign Ibjx84 = (Kcjx84 & Ytgx84);
	assign Kcjx84 = (~(S2jx84 & HRDATA[9]));
	assign K28x84 = (~(Rcjx84 & Ycjx84));
	assign Ycjx84 = (Ytgx84 & Wbjx84);
	assign Wbjx84 = (!S9jx84);
	assign S9jx84 = (Fdjx84 & Mdjx84);
	assign Fdjx84 = (~(Px0x84 | Kz0x84));
	assign Rcjx84 = (Tdjx84 & Aejx84);
	assign Aejx84 = (~(Kz0x84 & Hejx84));
	assign Hejx84 = (~(Oejx84 & Vejx84));
	assign Vejx84 = (~(Px0x84 & Glfx84));
	assign Tdjx84 = (~(S2jx84 & HRDATA[8]));
	assign E28x84 = (~(Cfjx84 & Jfjx84));
	assign Jfjx84 = (Px0x84 ? Oejx84 : Qfjx84);
	assign Oejx84 = (Ulfx84 & Xfjx84);
	assign Xfjx84 = (Mdjx84 | F6jx84);
	assign Cfjx84 = (Egjx84 & Ytgx84);
	assign Egjx84 = (~(S2jx84 & HRDATA[7]));
	assign Y18x84 = (~(Lgjx84 & Sgjx84));
	assign Sgjx84 = (Qfjx84 & Ytgx84);
	assign Ytgx84 = (~(W9ex84 & Zgjx84));
	assign Zgjx84 = (~(Ghjx84 & Nhjx84));
	assign Nhjx84 = (Uhjx84 & Bijx84);
	assign Bijx84 = (~(Iijx84 | Zt0x84));
	assign Iijx84 = (Tm0x84 ^ Pijx84);
	assign Uhjx84 = (Wijx84 & Dj0x84);
	assign Wijx84 = (~(Djjx84 ^ Oo0x84));
	assign Ghjx84 = (Kjjx84 & Rjjx84);
	assign Rjjx84 = (~(Yjjx84 ^ Yk0x84));
	assign Kjjx84 = (Fkjx84 & Mkjx84);
	assign Mkjx84 = (~(Tkjx84 ^ Jq0x84));
	assign Fkjx84 = (~(Aljx84 ^ Es0x84));
	assign Qfjx84 = (!Mdjx84);
	assign Mdjx84 = (Hljx84 & Dj0x84);
	assign Hljx84 = (~(Oljx84 | Uv0x84));
	assign Oljx84 = (!Vljx84);
	assign Lgjx84 = (Cmjx84 & Jmjx84);
	assign Jmjx84 = (~(S2jx84 & HRDATA[6]));
	assign Cmjx84 = (~(Uv0x84 & X1jx84));
	assign S18x84 = (~(Qmjx84 & Xmjx84));
	assign Xmjx84 = (~(S2jx84 & HRDATA[5]));
	assign Qmjx84 = (~(Zt0x84 & Enjx84));
	assign M18x84 = (~(Qrex84 & Lnjx84));
	assign Lnjx84 = (~(Snjx84 & Js3x84));
	assign Snjx84 = (Znjx84 & Gojx84);
	assign Gojx84 = (~(Ntex84 & HWDATA[25]));
	assign Znjx84 = (~(Nojx84 & Qcfx84));
	assign Qrex84 = (Uojx84 & Bpjx84);
	assign Bpjx84 = (~(Ipjx84 & Ppjx84));
	assign Ppjx84 = (Pu63a4[0] & Oo3x84);
	assign Ipjx84 = (Idhx84 & Pdhx84);
	assign Uojx84 = (~(Ntex84 & HWDATA[26]));
	assign Ntex84 = (Wpjx84 & In4w84);
	assign G18x84 = (Dqjx84 & Kqjx84);
	assign Kqjx84 = (Rqjx84 & Dgfx84);
	assign Dgfx84 = (~(HWDATA[2] & Wuex84));
	assign Rqjx84 = (~(Nmex84 & Yqjx84));
	assign Dqjx84 = (IRQ[2] & Frjx84);
	assign Frjx84 = (~(Pffx84 & Nefx84));
	assign Nefx84 = (~(Yqjx84 & Qcfx84));
	assign Pffx84 = (!Eu3x84);
	assign A18x84 = (Mrjx84 & Trjx84);
	assign Trjx84 = (Asjx84 & Cjfx84);
	assign Cjfx84 = (~(Wpjx84 & Szex84));
	assign Szex84 = (In4w84 & HWDATA[31]);
	assign Asjx84 = (Mpex84 | Cwgx84);
	assign Mrjx84 = (NMI & Hsjx84);
	assign Hsjx84 = (~(Vifx84 & Thfx84));
	assign Thfx84 = (Cwgx84 | Yoex84);
	assign Vifx84 = (!Ke63a4);
	assign U08x84 = (Osjx84 & Vsjx84);
	assign Vsjx84 = (~(Q5fx84 | Z6fx84));
	assign Z6fx84 = (HWDATA[1] & Wuex84);
	assign Q5fx84 = (N54x84 & E6fx84);
	assign E6fx84 = (~(Ctjx84 & Qcfx84));
	assign Osjx84 = (IRQ[1] & Jtjx84);
	assign Jtjx84 = (~(Nmex84 & Ctjx84));
	assign O08x84 = (~(Qtjx84 & Xtjx84));
	assign Xtjx84 = (Eujx84 & Lujx84);
	assign Lujx84 = (~(Kpdx84 & Qp63a4[9]));
	assign Eujx84 = (Sujx84 & Ypdx84);
	assign Sujx84 = (Igex84 | Bpcx84);
	assign Qtjx84 = (Zujx84 & Gvjx84);
	assign Gvjx84 = (~(Cr63a4[8] & Hrdx84));
	assign Zujx84 = (~(Tk63a4[8] & Ordx84));
	assign I08x84 = (~(Nvjx84 & Uvjx84));
	assign Uvjx84 = (Bwjx84 & Iwjx84);
	assign Iwjx84 = (~(Cr63a4[16] & Hrdx84));
	assign Bwjx84 = (Pwjx84 & Wwjx84);
	assign Wwjx84 = (Igex84 | Dxjx84);
	assign Pwjx84 = (~(Kpdx84 & Qp63a4[17]));
	assign Nvjx84 = (Jbgx84 & Kxjx84);
	assign Kxjx84 = (~(Tk63a4[16] & Ordx84));
	assign C08x84 = (~(Rxjx84 & Yxjx84));
	assign Yxjx84 = (Fyjx84 & Myjx84);
	assign Myjx84 = (~(Qp63a4[25] & Kpdx84));
	assign Fyjx84 = (Tyjx84 & Ypdx84);
	assign Tyjx84 = (Igex84 | Azjx84);
	assign Rxjx84 = (Hzjx84 & Ozjx84);
	assign Ozjx84 = (~(Cr63a4[24] & Hrdx84));
	assign Hzjx84 = (~(Tk63a4[24] & Ordx84));
	assign Wz7x84 = (Vzjx84 & C0kx84);
	assign C0kx84 = (~(D9fx84 | Tafx84));
	assign Tafx84 = (HWDATA[3] & Wuex84);
	assign Wuex84 = (C3hx84 & T8hx84);
	assign C3hx84 = (J0kx84 & In4w84);
	assign D9fx84 = (S54x84 & Q0kx84);
	assign Q0kx84 = (~(X0kx84 & Qcfx84));
	assign Vzjx84 = (IRQ[3] & E1kx84);
	assign E1kx84 = (Mpex84 | Y9fx84);
	assign Qz7x84 = (~(L1kx84 & S1kx84));
	assign S1kx84 = (Z1kx84 & G2kx84);
	assign G2kx84 = (~(Kpdx84 & Qp63a4[5]));
	assign Z1kx84 = (N2kx84 & Ypdx84);
	assign N2kx84 = (Igex84 | U2kx84);
	assign L1kx84 = (B3kx84 & I3kx84);
	assign I3kx84 = (~(Cr63a4[4] & Hrdx84));
	assign B3kx84 = (~(Tk63a4[4] & Ordx84));
	assign Kz7x84 = (~(P3kx84 & W3kx84));
	assign W3kx84 = (D4kx84 & K4kx84);
	assign K4kx84 = (~(Cr63a4[12] & Hrdx84));
	assign D4kx84 = (R4kx84 & Y4kx84);
	assign Y4kx84 = (Igex84 | F5kx84);
	assign R4kx84 = (~(Qp63a4[13] & Kpdx84));
	assign P3kx84 = (Wgex84 & M5kx84);
	assign M5kx84 = (~(Tk63a4[12] & Ordx84));
	assign Ez7x84 = (~(T5kx84 & A6kx84));
	assign A6kx84 = (H6kx84 & O6kx84);
	assign O6kx84 = (~(Cr63a4[20] & Hrdx84));
	assign H6kx84 = (V6kx84 & C7kx84);
	assign C7kx84 = (Igex84 | J7kx84);
	assign V6kx84 = (~(Qp63a4[21] & Kpdx84));
	assign T5kx84 = (Jbgx84 & Q7kx84);
	assign Q7kx84 = (~(Tk63a4[20] & Ordx84));
	assign Yy7x84 = (~(X7kx84 & E8kx84));
	assign E8kx84 = (L8kx84 & S8kx84);
	assign S8kx84 = (~(Qp63a4[2] & Kpdx84));
	assign L8kx84 = (Z8kx84 & Ypdx84);
	assign Z8kx84 = (Igex84 | G9kx84);
	assign X7kx84 = (N9kx84 & U9kx84);
	assign U9kx84 = (~(Cr63a4[1] & Hrdx84));
	assign N9kx84 = (~(V55w84 & Ordx84));
	assign Sy7x84 = (~(Bakx84 & Iakx84));
	assign Iakx84 = (Pakx84 & Wakx84);
	assign Wakx84 = (~(Cr63a4[9] & Hrdx84));
	assign Pakx84 = (Dbkx84 & Kbkx84);
	assign Kbkx84 = (Igex84 | Rbkx84);
	assign Dbkx84 = (~(Qp63a4[10] & Kpdx84));
	assign Bakx84 = (Wgex84 & Ybkx84);
	assign Ybkx84 = (~(Tk63a4[9] & Ordx84));
	assign My7x84 = (~(Fckx84 & Mckx84));
	assign Mckx84 = (Tckx84 & Adkx84);
	assign Adkx84 = (~(Cr63a4[17] & Hrdx84));
	assign Tckx84 = (Hdkx84 & Odkx84);
	assign Odkx84 = (Igex84 | Vdkx84);
	assign Hdkx84 = (~(Kpdx84 & Qp63a4[18]));
	assign Fckx84 = (Jbgx84 & Cekx84);
	assign Cekx84 = (~(Tk63a4[17] & Ordx84));
	assign Gy7x84 = (~(Jekx84 & Qekx84));
	assign Qekx84 = (Xekx84 & Efkx84);
	assign Efkx84 = (~(Qp63a4[26] & Kpdx84));
	assign Xekx84 = (Lfkx84 & Ypdx84);
	assign Lfkx84 = (Igex84 | Sfkx84);
	assign Jekx84 = (Zfkx84 & Ggkx84);
	assign Ggkx84 = (~(Cr63a4[25] & Hrdx84));
	assign Zfkx84 = (~(Tk63a4[25] & Ordx84));
	assign Ay7x84 = (~(Ngkx84 & Ugkx84));
	assign Ugkx84 = (~(Kf3x84 & Bhkx84));
	assign Bhkx84 = (~(Ihkx84 & Qcfx84));
	assign Qcfx84 = (!Yoex84);
	assign Ngkx84 = (Phkx84 | Zsex84);
	assign Zsex84 = (Whkx84 & Dikx84);
	assign Dikx84 = (~(Kikx84 & Hu2x84));
	assign Ux7x84 = (!Rikx84);
	assign Rikx84 = (X1jx84 ? Yikx84 : Glfx84);
	assign Yikx84 = (~(Fjkx84 & Ih0x84));
	assign Fjkx84 = (~(Mjkx84 | G8ex84));
	assign Glfx84 = (!F6jx84);
	assign Ox7x84 = (~(Tjkx84 & Akkx84));
	assign Akkx84 = (Hkkx84 & Okkx84);
	assign Okkx84 = (~(J6ex84 & HRDATA[30]));
	assign Hkkx84 = (Vkkx84 & Clkx84);
	assign Clkx84 = (~(K52x84 & E7ex84));
	assign Vkkx84 = (~(L7ex84 & HRDATA[14]));
	assign Tjkx84 = (Jlkx84 & Qlkx84);
	assign Qlkx84 = (~(Ka1x84 & G8ex84));
	assign Jlkx84 = (Xlkx84 | N8ex84);
	assign Ix7x84 = (~(Emkx84 & Lmkx84));
	assign Lmkx84 = (Smkx84 & Zmkx84);
	assign Zmkx84 = (~(HRDATA[28] & J6ex84));
	assign Smkx84 = (Gnkx84 & Nnkx84);
	assign Nnkx84 = (~(S12x84 & E7ex84));
	assign Gnkx84 = (~(HRDATA[12] & L7ex84));
	assign Emkx84 = (Unkx84 & Bokx84);
	assign Bokx84 = (~(S61x84 & G8ex84));
	assign Unkx84 = (Iokx84 | N8ex84);
	assign Cx7x84 = (~(Pokx84 & Wokx84));
	assign Wokx84 = (Dpkx84 & Kpkx84);
	assign Kpkx84 = (~(HRDATA[27] & J6ex84));
	assign Dpkx84 = (Rpkx84 & Ypkx84);
	assign Ypkx84 = (~(Wz1x84 & E7ex84));
	assign Rpkx84 = (~(HRDATA[11] & L7ex84));
	assign Pokx84 = (Fqkx84 & Mqkx84);
	assign Mqkx84 = (~(W41x84 & G8ex84));
	assign Fqkx84 = (Tqkx84 | N8ex84);
	assign Ww7x84 = (~(Arkx84 & Hrkx84));
	assign Hrkx84 = (Orkx84 & Vrkx84);
	assign Vrkx84 = (~(HRDATA[26] & J6ex84));
	assign Orkx84 = (Cskx84 & Jskx84);
	assign Jskx84 = (~(Ay1x84 & E7ex84));
	assign Cskx84 = (~(HRDATA[10] & L7ex84));
	assign Arkx84 = (Qskx84 & Xskx84);
	assign Xskx84 = (~(A31x84 & G8ex84));
	assign Qskx84 = (Tebx84 | N8ex84);
	assign Qw7x84 = (~(Etkx84 & Ltkx84));
	assign Ltkx84 = (Stkx84 & Ztkx84);
	assign Ztkx84 = (~(J6ex84 & HRDATA[25]));
	assign Stkx84 = (Gukx84 & Nukx84);
	assign Nukx84 = (~(Fw1x84 & E7ex84));
	assign Gukx84 = (~(L7ex84 & HRDATA[9]));
	assign Etkx84 = (Uukx84 & Bvkx84);
	assign Bvkx84 = (~(F11x84 & G8ex84));
	assign Uukx84 = (Wcbx84 | N8ex84);
	assign Kw7x84 = (~(Ivkx84 & Pvkx84));
	assign Pvkx84 = (Wvkx84 & Dwkx84);
	assign Dwkx84 = (~(J6ex84 & HRDATA[24]));
	assign Wvkx84 = (Kwkx84 & Rwkx84);
	assign Rwkx84 = (~(Ku1x84 & E7ex84));
	assign Kwkx84 = (~(L7ex84 & HRDATA[8]));
	assign Ivkx84 = (Ywkx84 & Fxkx84);
	assign Fxkx84 = (~(Kz0x84 & G8ex84));
	assign Ywkx84 = (Eobx84 | N8ex84);
	assign Ew7x84 = (~(Mxkx84 & Txkx84));
	assign Txkx84 = (Aykx84 & Hykx84);
	assign Hykx84 = (~(J6ex84 & HRDATA[23]));
	assign Aykx84 = (Oykx84 & Vykx84);
	assign Vykx84 = (~(Ps1x84 & E7ex84));
	assign Oykx84 = (~(L7ex84 & HRDATA[7]));
	assign Mxkx84 = (Czkx84 & Jzkx84);
	assign Jzkx84 = (~(Px0x84 & G8ex84));
	assign Czkx84 = (Qzkx84 | N8ex84);
	assign Yv7x84 = (~(Xzkx84 & E0lx84));
	assign E0lx84 = (L0lx84 & S0lx84);
	assign S0lx84 = (~(J6ex84 & HRDATA[22]));
	assign L0lx84 = (Z0lx84 & G1lx84);
	assign G1lx84 = (~(Uq1x84 & E7ex84));
	assign Z0lx84 = (~(L7ex84 & HRDATA[6]));
	assign Xzkx84 = (N1lx84 & U1lx84);
	assign U1lx84 = (~(Uv0x84 & G8ex84));
	assign N1lx84 = (Jfcx84 | N8ex84);
	assign Sv7x84 = (~(B2lx84 & I2lx84));
	assign I2lx84 = (P2lx84 & W2lx84);
	assign W2lx84 = (~(HRDATA[21] & J6ex84));
	assign P2lx84 = (D3lx84 & K3lx84);
	assign K3lx84 = (~(Zo1x84 & E7ex84));
	assign D3lx84 = (~(HRDATA[5] & L7ex84));
	assign B2lx84 = (R3lx84 & Y3lx84);
	assign Y3lx84 = (~(G8ex84 & Zt0x84));
	assign R3lx84 = (Iicx84 | N8ex84);
	assign Mv7x84 = (~(F4lx84 & M4lx84));
	assign M4lx84 = (T4lx84 & A5lx84);
	assign A5lx84 = (~(HRDATA[20] & J6ex84));
	assign T4lx84 = (H5lx84 & O5lx84);
	assign O5lx84 = (~(En1x84 & E7ex84));
	assign H5lx84 = (~(HRDATA[4] & L7ex84));
	assign F4lx84 = (V5lx84 & C6lx84);
	assign C6lx84 = (~(Es0x84 & G8ex84));
	assign V5lx84 = (Jmcx84 | N8ex84);
	assign Gv7x84 = (~(Puex84 & J6lx84));
	assign J6lx84 = (~(Cc3x84 & Q6lx84));
	assign Q6lx84 = (~(X6lx84 & Nj63a4[0]));
	assign X6lx84 = (~(Yoex84 | E7lx84));
	assign Yoex84 = (~(L7lx84 & Zo2x84));
	assign L7lx84 = (~(T7bx84 | N4ix84));
	assign Puex84 = (S7lx84 & Z7lx84);
	assign Z7lx84 = (Whkx84 | Ssex84);
	assign Whkx84 = (~(G8lx84 & N8lx84));
	assign N8lx84 = (~(S1dx84 | N4ix84));
	assign G8lx84 = (U8lx84 & B9lx84);
	assign S7lx84 = (I9lx84 & P9lx84);
	assign P9lx84 = (~(W9lx84 & Dalx84));
	assign Dalx84 = (Kalx84 & Ralx84);
	assign Kalx84 = (Hscx84 | E7lx84);
	assign W9lx84 = (~(H6dx84 | Ambx84));
	assign I9lx84 = (~(Yalx84 & Vvgx84));
	assign Yalx84 = (~(Fblx84 & Mblx84));
	assign Fblx84 = (Tblx84 & Aclx84);
	assign Aclx84 = (~(Hclx84 & D53x84));
	assign Hclx84 = (~(Ambx84 | Ralx84));
	assign Tblx84 = (~(Oclx84 & Tsix84));
	assign Av7x84 = (Vclx84 ? Lmdx84 : SLEEPHOLDREQn);
	assign Vclx84 = (Cdlx84 & Jdlx84);
	assign Jdlx84 = (~(Qdlx84 & Xdlx84));
	assign Xdlx84 = (~(Eelx84 & Lelx84));
	assign Cdlx84 = (~(SLEEPHOLDREQn & HREADY));
	assign Uu7x84 = (~(Selx84 & Zelx84));
	assign Zelx84 = (Gflx84 & Nflx84);
	assign Nflx84 = (~(HRDATA[19] & J6ex84));
	assign Gflx84 = (Uflx84 & Bglx84);
	assign Bglx84 = (~(Jl1x84 & E7ex84));
	assign Uflx84 = (~(HRDATA[3] & L7ex84));
	assign Selx84 = (Iglx84 & Pglx84);
	assign Pglx84 = (~(Jq0x84 & G8ex84));
	assign Iglx84 = (Rufx84 | N8ex84);
	assign Ou7x84 = (~(Wglx84 & Dhlx84));
	assign Dhlx84 = (Khlx84 & Rhlx84);
	assign Rhlx84 = (~(Czdx84 & Nj63a4[2]));
	assign Khlx84 = (~(Jzdx84 & HADDR[2]));
	assign Wglx84 = (Yhlx84 & Filx84);
	assign Filx84 = (~(E0ex84 & V55w84));
	assign Yhlx84 = (~(S09w84 & L0ex84));
	assign Iu7x84 = (~(Milx84 & Tilx84));
	assign Tilx84 = (Ajlx84 & Hjlx84);
	assign Hjlx84 = (~(HRDATA[18] & J6ex84));
	assign Ajlx84 = (Ojlx84 & Vjlx84);
	assign Vjlx84 = (~(Oj1x84 & E7ex84));
	assign Ojlx84 = (~(HRDATA[2] & L7ex84));
	assign Milx84 = (Cklx84 & Jklx84);
	assign Jklx84 = (~(Oo0x84 & G8ex84));
	assign Cklx84 = (Qklx84 | N8ex84);
	assign Cu7x84 = (~(Xklx84 & Ellx84));
	assign Ellx84 = (Lllx84 & Sllx84);
	assign Sllx84 = (~(J6ex84 & HRDATA[17]));
	assign J6ex84 = (Zllx84 & Gmlx84);
	assign Lllx84 = (Nmlx84 & Umlx84);
	assign Umlx84 = (~(Th1x84 & E7ex84));
	assign E7ex84 = (Bnlx84 & N8ex84);
	assign Bnlx84 = (Inlx84 & Wmfx84);
	assign Inlx84 = (~(Prax84 & Pnlx84));
	assign Pnlx84 = (Bzgx84 | Ih0x84);
	assign Nmlx84 = (~(L7ex84 & HRDATA[1]));
	assign L7ex84 = (Zllx84 & Wnlx84);
	assign Wnlx84 = (~(Wmfx84 | Gmlx84));
	assign Gmlx84 = (Tk63a4[0] & Gpbx84);
	assign Wmfx84 = (!Ya2x84);
	assign Zllx84 = (~(Nlfx84 | Dolx84));
	assign Xklx84 = (Kolx84 & Rolx84);
	assign Rolx84 = (~(Tm0x84 & G8ex84));
	assign G8ex84 = (Ih0x84 & N8ex84);
	assign Kolx84 = (Yufx84 | N8ex84);
	assign N8ex84 = (!Dolx84);
	assign Dolx84 = (~(Yolx84 & Fplx84));
	assign Fplx84 = (Mplx84 & Tplx84);
	assign Mplx84 = (~(Aqlx84 | LOCKUP));
	assign Yolx84 = (O2hx84 & Hqlx84);
	assign Hqlx84 = (~(Oqlx84 & Qwgx84));
	assign Oqlx84 = (~(Vqlx84 & Crlx84));
	assign Vqlx84 = (Prax84 & Jrlx84);
	assign Wt7x84 = (Csdx84 ? Km63a4[3] : Qrlx84);
	assign Qrlx84 = (~(Ztdx84 & Xrlx84));
	assign Xrlx84 = (~(G36w84 & Eslx84));
	assign Eslx84 = (~(Saix84 & Lslx84));
	assign Lslx84 = (~(Sslx84 & I86w84));
	assign Qt7x84 = (Csdx84 ? Km63a4[2] : Zslx84);
	assign Zslx84 = (~(Gtlx84 & Ntlx84));
	assign Ntlx84 = (Utlx84 & Bulx84);
	assign Bulx84 = (~(Wz5w84 & Ltdx84));
	assign Utlx84 = (~(Uu5w84 & Stdx84));
	assign Gtlx84 = (Ztdx84 & Iulx84);
	assign Iulx84 = (~(I86w84 & Nudx84));
	assign Ztdx84 = (Pulx84 & Wulx84);
	assign Wulx84 = (Dvlx84 & Kvlx84);
	assign Kvlx84 = (~(Rvlx84 | Gwix84));
	assign Dvlx84 = (Yvlx84 & Zrfx84);
	assign Zrfx84 = (J13x84 | E8dx84);
	assign Yvlx84 = (~(Zg6w84 & Fwlx84));
	assign Fwlx84 = (~(Leex84 ^ Ub6w84));
	assign Pulx84 = (Mwlx84 & Twlx84);
	assign Mwlx84 = (Axlx84 & Hxlx84);
	assign Hxlx84 = (~(Oxlx84 & Wcbx84));
	assign Axlx84 = (Rufx84 | Ambx84);
	assign Kt7x84 = (Csdx84 ? Km63a4[1] : Vxlx84);
	assign Csdx84 = (~(HREADY & Cylx84));
	assign Cylx84 = (~(Jylx84 & Qylx84));
	assign Qylx84 = (Xylx84 & Ezlx84);
	assign Ezlx84 = (~(Lzlx84 & Szlx84));
	assign Szlx84 = (~(Zzlx84 & G0mx84));
	assign G0mx84 = (N0mx84 | Gpbx84);
	assign Xylx84 = (U0mx84 & Mpex84);
	assign Mpex84 = (!Nmex84);
	assign Nmex84 = (Afix84 & Pqbx84);
	assign U0mx84 = (~(Nzfx84 & B1mx84));
	assign B1mx84 = (~(B0gx84 & I1mx84));
	assign I1mx84 = (P1mx84 | Gz4w84);
	assign Jylx84 = (W1mx84 & D2mx84);
	assign W1mx84 = (K2mx84 & R2mx84);
	assign R2mx84 = (~(Y2mx84 & F3mx84));
	assign Y2mx84 = (~(M3mx84 & T3mx84));
	assign T3mx84 = (A4mx84 & H4mx84);
	assign H4mx84 = (~(L2cx84 & O4mx84));
	assign O4mx84 = (Xlkx84 | Mcdx84);
	assign A4mx84 = (V4mx84 & C5mx84);
	assign V4mx84 = (~(J5mx84 & Q5mx84));
	assign Q5mx84 = (G36w84 | Ba6w84);
	assign M3mx84 = (X5mx84 & E6mx84);
	assign E6mx84 = (~(L6mx84 & S6mx84));
	assign X5mx84 = (~(V1ix84 & Z6mx84));
	assign K2mx84 = (Mzbx84 | Dybx84);
	assign Vxlx84 = (~(G7mx84 & N7mx84));
	assign N7mx84 = (U7mx84 & B8mx84);
	assign B8mx84 = (~(Ey5w84 & Ltdx84));
	assign Ltdx84 = (~(I8mx84 & P8mx84));
	assign P8mx84 = (~(W8mx84 & D9mx84));
	assign I8mx84 = (~(K9mx84 & Ambx84));
	assign K9mx84 = (Nd6w84 ? Y9mx84 : R9mx84);
	assign Y9mx84 = (~(Famx84 & Ouhx84));
	assign Famx84 = (~(Mamx84 & Q66w84));
	assign Mamx84 = (Oxlx84 & E8dx84);
	assign R9mx84 = (Tamx84 & Xlkx84);
	assign U7mx84 = (~(Ct5w84 & Stdx84));
	assign Stdx84 = (Sslx84 | Abmx84);
	assign Abmx84 = (Hbmx84 & Rufx84);
	assign G7mx84 = (Twlx84 & Obmx84);
	assign Obmx84 = (~(Q66w84 & Nudx84));
	assign Nudx84 = (~(Vbmx84 & Ccmx84));
	assign Ccmx84 = (~(Jcmx84 & Nd6w84));
	assign Jcmx84 = (~(Qcmx84 | Xcmx84));
	assign Vbmx84 = (~(Edmx84 & Ambx84));
	assign Twlx84 = (Ldmx84 & Sdmx84);
	assign Sdmx84 = (~(Zdmx84 & Sslx84));
	assign Sslx84 = (Gemx84 & Nemx84);
	assign Nemx84 = (~(Ub6w84 | Nd6w84));
	assign Gemx84 = (Uemx84 & D9mx84);
	assign Zdmx84 = (Bfmx84 & Ifmx84);
	assign Ldmx84 = (Pfmx84 & Wfmx84);
	assign Wfmx84 = (~(Ambx84 & Dgmx84));
	assign Dgmx84 = (~(Kgmx84 & Rgmx84));
	assign Rgmx84 = (~(Ygmx84 & Lzlx84));
	assign Ygmx84 = (Nd6w84 & Tamx84);
	assign Kgmx84 = (~(Fhmx84 & Oxlx84));
	assign Pfmx84 = (~(Mhmx84 & Thmx84));
	assign Thmx84 = (~(Kr5w84 | Ct5w84));
	assign Mhmx84 = (~(Rufx84 | Saix84));
	assign Et7x84 = (Himx84 ? Aimx84 : O75w84);
	assign Aimx84 = (~(Oimx84 & Vimx84));
	assign Vimx84 = (Cjmx84 & Jjmx84);
	assign Jjmx84 = (Qjmx84 & Niix84);
	assign Qjmx84 = (~(Xjmx84 & Ekmx84));
	assign Xjmx84 = (~(Lkmx84 & Skmx84));
	assign Skmx84 = (Kkbx84 | Iv6w84);
	assign Lkmx84 = (Zkmx84 & Glmx84);
	assign Glmx84 = (~(Nlmx84 & Kjcx84));
	assign Zkmx84 = (Sgcx84 | Ulmx84);
	assign Cjmx84 = (Bmmx84 & Immx84);
	assign Immx84 = (~(Mw5w84 & Pmmx84));
	assign Bmmx84 = (Wmmx84 | Dnmx84);
	assign Oimx84 = (Knmx84 & Rnmx84);
	assign Knmx84 = (Ynmx84 & Fomx84);
	assign Fomx84 = (~(Momx84 & Kr5w84));
	assign Ynmx84 = (Cgix84 | Jfcx84);
	assign Ys7x84 = (Gqhx84 ? Tomx84 : Ln6w84);
	assign Tomx84 = (~(Apmx84 & Hpmx84));
	assign Hpmx84 = (Opmx84 & Vpmx84);
	assign Vpmx84 = (Cqmx84 & Jqmx84);
	assign Jqmx84 = (~(Qqmx84 & Xqmx84));
	assign Cqmx84 = (Ermx84 & Lrmx84);
	assign Lrmx84 = (~(Srmx84 & Cvhx84));
	assign Srmx84 = (Zrmx84 | Gsmx84);
	assign Gsmx84 = (~(Nsmx84 | Usmx84));
	assign Ermx84 = (~(Btmx84 & F7ix84));
	assign Btmx84 = (~(Itmx84 ^ I3dx84));
	assign Opmx84 = (Ptmx84 & Wtmx84);
	assign Wtmx84 = (~(Dumx84 & Uu5w84));
	assign Ptmx84 = (Kumx84 & Rumx84);
	assign Rumx84 = (~(Q66w84 & Yumx84));
	assign Kumx84 = (~(Lwhx84 & Jq0x84));
	assign Apmx84 = (Fvmx84 & Mvmx84);
	assign Mvmx84 = (Tvmx84 & Awmx84);
	assign Awmx84 = (~(W05w84 & Hwmx84));
	assign Tvmx84 = (Owmx84 & Vwmx84);
	assign Vwmx84 = (Rufx84 | Byhx84);
	assign Owmx84 = (Lncx84 | Eobx84);
	assign Fvmx84 = (Uiix84 & Cxmx84);
	assign Cxmx84 = (Jxmx84 | Qxmx84);
	assign Uiix84 = (Xxmx84 & Eymx84);
	assign Eymx84 = (~(Lymx84 & W05w84));
	assign Lymx84 = (F7bx84 & Yqcx84);
	assign Xxmx84 = (~(Symx84 | Zymx84));
	assign Ss7x84 = (~(Gzmx84 & Nzmx84));
	assign Nzmx84 = (~(Wl6w84 & Uzmx84));
	assign Uzmx84 = (~(Gqhx84 & B0nx84));
	assign B0nx84 = (Iyhx84 | I0nx84);
	assign Gzmx84 = (~(Gqhx84 & P0nx84));
	assign P0nx84 = (~(W0nx84 & D1nx84));
	assign D1nx84 = (K1nx84 & R1nx84);
	assign R1nx84 = (Y1nx84 & F2nx84);
	assign F2nx84 = (~(M2nx84 & I0nx84));
	assign M2nx84 = (~(Iyhx84 | Wl6w84));
	assign Iyhx84 = (!F7ix84);
	assign Y1nx84 = (~(T2nx84 & Cvhx84));
	assign T2nx84 = (~(Nsmx84 ^ A3nx84));
	assign A3nx84 = (~(Zrmx84 | Usmx84));
	assign Usmx84 = (H3nx84 & O3nx84);
	assign O3nx84 = (V3nx84 & C4nx84);
	assign H3nx84 = (J4nx84 & Q4nx84);
	assign Q4nx84 = (~(X4nx84 & E5nx84));
	assign Zrmx84 = (L5nx84 & X4nx84);
	assign L5nx84 = (E5nx84 & S5nx84);
	assign S5nx84 = (~(J4nx84 & V3nx84));
	assign V3nx84 = (Z5nx84 | G6nx84);
	assign J4nx84 = (N6nx84 & U6nx84);
	assign N6nx84 = (B7nx84 | I7nx84);
	assign K1nx84 = (P7nx84 & W7nx84);
	assign W7nx84 = (~(Lwhx84 & Oo0x84));
	assign P7nx84 = (~(Y46w84 & Swhx84));
	assign W0nx84 = (D8nx84 & K8nx84);
	assign K8nx84 = (R8nx84 & Y8nx84);
	assign Y8nx84 = (~(Dumx84 & Ct5w84));
	assign R8nx84 = (Qklx84 | Byhx84);
	assign D8nx84 = (Dzhx84 & F9nx84);
	assign F9nx84 = (Lncx84 | Qzkx84);
	assign Ms7x84 = (~(M9nx84 & T9nx84));
	assign T9nx84 = (~(Aanx84 & F7ix84));
	assign M9nx84 = (Gqhx84 ? Oanx84 : Hanx84);
	assign Gqhx84 = (HREADY & Vanx84);
	assign Vanx84 = (~(Cbnx84 & Jbnx84));
	assign Jbnx84 = (Qbnx84 & Xbnx84);
	assign Xbnx84 = (Ecnx84 & Lcnx84);
	assign Qbnx84 = (Scnx84 & Zcnx84);
	assign Zcnx84 = (~(Gdnx84 & Ndnx84));
	assign Ndnx84 = (~(Evix84 | Gz4w84));
	assign Gdnx84 = (Nacx84 & Undx84);
	assign Scnx84 = (~(Udnx84 & Benx84));
	assign Udnx84 = (~(Tebx84 | W05w84));
	assign Cbnx84 = (Ienx84 & Penx84);
	assign Penx84 = (Wenx84 & Dfnx84);
	assign Dfnx84 = (~(Kfnx84 & Rfnx84));
	assign Kfnx84 = (~(Tsix84 | Vx2x84));
	assign Wenx84 = (~(Yfnx84 & N4ix84));
	assign Yfnx84 = (~(Fthx84 | Wqbx84));
	assign Ienx84 = (Z3ix84 & Fgnx84);
	assign Fgnx84 = (~(A7cx84 & Mgnx84));
	assign Z3ix84 = (Tgnx84 & Ahnx84);
	assign Ahnx84 = (Hhnx84 & Ohnx84);
	assign Ohnx84 = (Vhnx84 & Cinx84);
	assign Cinx84 = (~(Jinx84 & Lzlx84));
	assign Jinx84 = (Gz4w84 & Qinx84);
	assign Qinx84 = (~(Xlkx84 & Xinx84));
	assign Xinx84 = (Y46w84 | Q66w84);
	assign Vhnx84 = (~(Ejnx84 | Ljnx84));
	assign Hhnx84 = (Sjnx84 & Zjnx84);
	assign Zjnx84 = (~(Nzfx84 & Gknx84));
	assign Sjnx84 = (Nknx84 & Uknx84);
	assign Uknx84 = (~(Blnx84 & Ilnx84));
	assign Blnx84 = (Plnx84 & Rufx84);
	assign Nknx84 = (~(Wlnx84 & Dmnx84));
	assign Dmnx84 = (~(Y4dx84 & Kmnx84));
	assign Kmnx84 = (Rmnx84 | Jxmx84);
	assign Tgnx84 = (Ymnx84 & Fnnx84);
	assign Fnnx84 = (Mnnx84 & Tnnx84);
	assign Mnnx84 = (Aonx84 & Honx84);
	assign Honx84 = (~(Oonx84 & F3mx84));
	assign Oonx84 = (~(Vonx84 & Cpnx84));
	assign Cpnx84 = (~(Jpnx84 & Xlkx84));
	assign Vonx84 = (Qpnx84 & C5mx84);
	assign Qpnx84 = (~(L2cx84 & Xpnx84));
	assign Xpnx84 = (~(Eqnx84 & Lqnx84));
	assign Lqnx84 = (~(Sqnx84 & Zqnx84));
	assign Zqnx84 = (~(Qzkx84 | Ba6w84));
	assign Sqnx84 = (~(Eobx84 | Z6mx84));
	assign Eqnx84 = (~(Grnx84 & Nrnx84));
	assign Ymnx84 = (Urnx84 & Bsnx84);
	assign Oanx84 = (Isnx84 & Psnx84);
	assign Psnx84 = (Wsnx84 & Dtnx84);
	assign Dtnx84 = (Ktnx84 & Rtnx84);
	assign Rtnx84 = (~(Ytnx84 & Funx84));
	assign Funx84 = (~(Munx84 & Tunx84));
	assign Tunx84 = (~(Qvhx84 & Jvhx84));
	assign Munx84 = (~(X4nx84 ^ E5nx84));
	assign Ytnx84 = (Nsmx84 & Cvhx84);
	assign Cvhx84 = (~(Avnx84 & Hvnx84));
	assign Hvnx84 = (~(Ovnx84 & I86w84));
	assign Avnx84 = (~(Shix84 & Edmx84));
	assign Nsmx84 = (~(Vvnx84 & Qvhx84));
	assign Qvhx84 = (~(Eobx84 | Iokx84));
	assign Vvnx84 = (E5nx84 & Jvhx84);
	assign Jvhx84 = (~(Cwnx84 | X4nx84));
	assign X4nx84 = (G36w84 & Jwnx84);
	assign Jwnx84 = (Jfcx84 ^ Qwnx84);
	assign Cwnx84 = (Xwnx84 & Qzkx84);
	assign Xwnx84 = (~(Qwnx84 ^ Jfcx84));
	assign E5nx84 = (Exnx84 & C4nx84);
	assign C4nx84 = (Lxnx84 | I7nx84);
	assign Exnx84 = (~(Sxnx84 & Lxnx84));
	assign Lxnx84 = (Qwnx84 | Jfcx84);
	assign Qwnx84 = (~(Zxnx84 & B7nx84));
	assign Zxnx84 = (~(Gynx84 & Iicx84));
	assign Sxnx84 = (~(I7nx84 ^ B7nx84));
	assign B7nx84 = (Iicx84 | Gynx84);
	assign Gynx84 = (Nynx84 ^ Jmcx84);
	assign I7nx84 = (~(Uynx84 & U6nx84));
	assign U6nx84 = (~(Bznx84 & Nynx84));
	assign Bznx84 = (~(Jmcx84 | G6nx84));
	assign Uynx84 = (~(Iznx84 & Pznx84));
	assign Pznx84 = (~(Nynx84 & Ey5w84));
	assign Nynx84 = (Z5nx84 & Wznx84);
	assign Wznx84 = (~(D0ox84 & Rufx84));
	assign Iznx84 = (~(G6nx84 ^ Z5nx84));
	assign Z5nx84 = (D0ox84 | Rufx84);
	assign D0ox84 = (K0ox84 | R0ox84);
	assign K0ox84 = (Y0ox84 & Qklx84);
	assign G6nx84 = (~(F1ox84 | R0ox84));
	assign R0ox84 = (~(Qklx84 | Y0ox84));
	assign Y0ox84 = (~(Kr5w84 ^ Ct5w84));
	assign Ktnx84 = (~(Lwhx84 & Tm0x84));
	assign Lwhx84 = (Dj0x84 & M1ox84);
	assign M1ox84 = (~(T1ox84 & Meix84));
	assign Meix84 = (Jxmx84 | A2ox84);
	assign T1ox84 = (H2ox84 & O2ox84);
	assign H2ox84 = (Yqcx84 | V2ox84);
	assign Wsnx84 = (C3ox84 & J3ox84);
	assign J3ox84 = (~(G36w84 & Swhx84));
	assign Swhx84 = (Yumx84 | Xqmx84);
	assign Yumx84 = (~(Bcix84 & Q3ox84));
	assign Q3ox84 = (~(Pcix84 & Huhx84));
	assign C3ox84 = (~(Dumx84 & Kr5w84));
	assign Dumx84 = (Fhmx84 & X3ox84);
	assign X3ox84 = (~(Cgix84 & E4ox84));
	assign E4ox84 = (L4ox84 | Gpbx84);
	assign Isnx84 = (S4ox84 & Z4ox84);
	assign Z4ox84 = (G5ox84 & N5ox84);
	assign N5ox84 = (Yufx84 | Byhx84);
	assign Byhx84 = (U5ox84 & B6ox84);
	assign B6ox84 = (I6ox84 & P6ox84);
	assign P6ox84 = (~(W6ox84 & D7ox84));
	assign D7ox84 = (~(Ouhx84 | Zg6w84));
	assign W6ox84 = (V1ix84 & Ba6w84);
	assign I6ox84 = (~(Kikx84 & E8dx84));
	assign U5ox84 = (Zhix84 & K7ox84);
	assign K7ox84 = (Cfcx84 | I86w84);
	assign Zhix84 = (R7ox84 & Y7ox84);
	assign Y7ox84 = (~(Pcix84 & F8ox84));
	assign Yufx84 = (!Ct5w84);
	assign G5ox84 = (~(M8ox84 & F7ix84));
	assign F7ix84 = (~(T8ox84 & A9ox84));
	assign A9ox84 = (H9ox84 & O9ox84);
	assign O9ox84 = (V9ox84 & Erfx84);
	assign Erfx84 = (~(Caox84 & J13x84));
	assign Caox84 = (~(Tq2x84 | Ns2x84));
	assign H9ox84 = (Jaox84 & Qaox84);
	assign Qaox84 = (~(Mlbx84 & Xaox84));
	assign Xaox84 = (~(Ebox84 & Lbox84));
	assign Lbox84 = (Sbox84 | Cuix84);
	assign Jaox84 = (Saix84 | Zbox84);
	assign T8ox84 = (Gcox84 & Ncox84);
	assign Ncox84 = (Ucox84 | Bdox84);
	assign Gcox84 = (Idox84 & Pdox84);
	assign Pdox84 = (~(U8lx84 & Wdox84));
	assign Idox84 = (~(Rzhx84 & Deox84));
	assign S4ox84 = (Dzhx84 & Keox84);
	assign Keox84 = (Lncx84 | Jfcx84);
	assign Dzhx84 = (Reox84 & Yeox84);
	assign Yeox84 = (V2ox84 | Tq2x84);
	assign Reox84 = (~(Ffox84 & Uu5w84));
	assign Gs7x84 = (Himx84 ? Mfox84 : H95w84);
	assign Mfox84 = (~(Tfox84 & Agox84));
	assign Agox84 = (Hgox84 & Ogox84);
	assign Ogox84 = (Wmmx84 | Kkbx84);
	assign Hgox84 = (Vgox84 & Chox84);
	assign Chox84 = (~(Jhox84 & Ekmx84));
	assign Jhox84 = (~(Kjcx84 & Qhox84));
	assign Qhox84 = (~(Xhox84 & Vfbx84));
	assign Vgox84 = (~(Ey5w84 & Pmmx84));
	assign Tfox84 = (Eiox84 & Rnmx84);
	assign Rnmx84 = (Liox84 & Siox84);
	assign Siox84 = (~(Ziox84 & Gjox84));
	assign Ziox84 = (Ekmx84 & C9ix84);
	assign C9ix84 = (!Njox84);
	assign Eiox84 = (Ujox84 & Bkox84);
	assign Bkox84 = (~(Momx84 & Ct5w84));
	assign Ujox84 = (Cgix84 | Qzkx84);
	assign As7x84 = (Himx84 ? Ikox84 : Ab5w84);
	assign Ikox84 = (~(Pkox84 & Wkox84));
	assign Wkox84 = (Dlox84 & Klox84);
	assign Klox84 = (Rlox84 & Niix84);
	assign Rlox84 = (~(Wz5w84 & Pmmx84));
	assign Pmmx84 = (~(Zzlx84 & Ylox84));
	assign Ylox84 = (E2cx84 | Tebx84);
	assign Dlox84 = (Fmox84 & Mmox84);
	assign Mmox84 = (~(Njox84 & Ekmx84));
	assign Fmox84 = (Wmmx84 | Tmox84);
	assign Pkox84 = (Anox84 & Liox84);
	assign Anox84 = (Hnox84 & Onox84);
	assign Onox84 = (~(Momx84 & Uu5w84));
	assign Hnox84 = (Eobx84 | Cgix84);
	assign Ur7x84 = (Himx84 ? Vnox84 : Tc5w84);
	assign Himx84 = (~(Coox84 & Joox84));
	assign Joox84 = (~(Qoox84 & Xoox84));
	assign Xoox84 = (~(Epox84 & Lpox84));
	assign Lpox84 = (~(Frcx84 & Spox84));
	assign Epox84 = (Zpox84 & Gqox84);
	assign Zpox84 = (~(Nqox84 & N4ix84));
	assign Nqox84 = (~(Fthx84 | Jnix84));
	assign Coox84 = (~(HREADY & Uqox84));
	assign Uqox84 = (~(Brox84 & Irox84));
	assign Irox84 = (Prox84 & Wrox84);
	assign Wrox84 = (Dsox84 & Ksox84);
	assign Ksox84 = (~(Rsox84 & Lfdx84));
	assign Rsox84 = (Ysox84 & Iicx84);
	assign Dsox84 = (Ftox84 & Mtox84);
	assign Ftox84 = (~(Ttox84 & Auox84));
	assign Ttox84 = (Huox84 & Mw5w84);
	assign Prox84 = (Ouox84 & Vuox84);
	assign Vuox84 = (~(Cvox84 & Yrbx84));
	assign Cvox84 = (Nwix84 & Iqbx84);
	assign Ouox84 = (Jvox84 & Qvox84);
	assign Qvox84 = (~(Xvox84 & Xqmx84));
	assign Xvox84 = (Ewox84 & F3mx84);
	assign Ewox84 = (~(Xlkx84 & Lwox84));
	assign Lwox84 = (Tqkx84 | I86w84);
	assign Jvox84 = (~(Swox84 & Jpnx84));
	assign Swox84 = (Uemx84 & E8dx84);
	assign Brox84 = (Zwox84 & Gxox84);
	assign Gxox84 = (Nxox84 & Uxox84);
	assign Uxox84 = (~(Mlbx84 & Byox84));
	assign Byox84 = (~(Iyox84 & Pyox84));
	assign Pyox84 = (~(Frcx84 & Fn2x84));
	assign Iyox84 = (~(Wyox84 | Dzox84));
	assign Nxox84 = (Kzox84 & Rzox84);
	assign Rzox84 = (~(Yzox84 & Gwix84));
	assign Yzox84 = (~(Fthx84 | S1dx84));
	assign Kzox84 = (~(Rzhx84 & F0px84));
	assign F0px84 = (M0px84 | T0px84);
	assign Zwox84 = (A1px84 & H1px84);
	assign H1px84 = (Saix84 | O1px84);
	assign Vnox84 = (~(V1px84 & C2px84));
	assign C2px84 = (J2px84 & Q2px84);
	assign Q2px84 = (~(X2px84 & Ekmx84));
	assign Ekmx84 = (~(E3px84 & L3px84));
	assign L3px84 = (S3px84 & Ambx84);
	assign S3px84 = (~(Z3px84 & F2gx84));
	assign E3px84 = (G4px84 & N4px84);
	assign N4px84 = (U4px84 | Hu2x84);
	assign G4px84 = (A0cx84 | Bw2x84);
	assign X2px84 = (~(Akdx84 & B5px84));
	assign B5px84 = (~(I5px84 & Njox84));
	assign I5px84 = (~(D8gx84 | Ambx84));
	assign J2px84 = (P5px84 & Niix84);
	assign P5px84 = (~(W5px84 & I86w84));
	assign W5px84 = (O16w84 & D6px84);
	assign D6px84 = (L2cx84 | F8ox84);
	assign V1px84 = (K6px84 & Liox84);
	assign Liox84 = (R6px84 & Y6px84);
	assign Y6px84 = (Jxmx84 | Pz2x84);
	assign R6px84 = (Ecnx84 & Mzbx84);
	assign Ecnx84 = (Ambx84 | Dybx84);
	assign K6px84 = (F7px84 & M7px84);
	assign M7px84 = (Wmmx84 | T7px84);
	assign Wmmx84 = (~(Pxbx84 & A8px84));
	assign A8px84 = (H8px84 | O8px84);
	assign F7px84 = (~(Momx84 & Mw5w84));
	assign Or7x84 = (V8px84 ? C4uw84 : Wdhx84);
	assign Ir7x84 = (V8px84 ? X5uw84 : L5gx84);
	assign Cr7x84 = (V8px84 ? S7uw84 : F9gx84);
	assign Wq7x84 = (V8px84 ? Eavw84 : Xbgx84);
	assign Qq7x84 = (V8px84 ? Cnvw84 : Q4gx84);
	assign Kq7x84 = (V8px84 ? Yovw84 : E5gx84);
	assign Eq7x84 = (C9px84 ? Suqw84 : Wdhx84);
	assign Yp7x84 = (C9px84 ? Nwqw84 : L5gx84);
	assign Sp7x84 = (C9px84 ? Iyqw84 : F9gx84);
	assign Mp7x84 = (C9px84 ? U0sw84 : Xbgx84);
	assign Gp7x84 = (C9px84 ? Sdsw84 : Q4gx84);
	assign Ap7x84 = (C9px84 ? Ofsw84 : E5gx84);
	assign Uo7x84 = (J9px84 ? A8pw84 : Wdhx84);
	assign Oo7x84 = (J9px84 ? V9pw84 : L5gx84);
	assign Io7x84 = (J9px84 ? Qbpw84 : F9gx84);
	assign Co7x84 = (J9px84 ? Ceqw84 : Xbgx84);
	assign Wn7x84 = (J9px84 ? Arqw84 : Q4gx84);
	assign Qn7x84 = (J9px84 ? Wsqw84 : E5gx84);
	assign Kn7x84 = (Q9px84 ? Ilnw84 : Wdhx84);
	assign En7x84 = (Q9px84 ? Dnnw84 : L5gx84);
	assign Ym7x84 = (Q9px84 ? Yonw84 : F9gx84);
	assign Sm7x84 = (Q9px84 ? Krow84 : Xbgx84);
	assign Mm7x84 = (Q9px84 ? I4pw84 : Q4gx84);
	assign Gm7x84 = (Q9px84 ? E6pw84 : E5gx84);
	assign Am7x84 = (X9px84 ? Qylw84 : Wdhx84);
	assign Ul7x84 = (X9px84 ? L0mw84 : L5gx84);
	assign Ol7x84 = (X9px84 ? G2mw84 : F9gx84);
	assign Il7x84 = (X9px84 ? S4nw84 : Xbgx84);
	assign Cl7x84 = (X9px84 ? Qhnw84 : Q4gx84);
	assign Wk7x84 = (X9px84 ? Mjnw84 : E5gx84);
	assign Qk7x84 = (Eapx84 ? Ybkw84 : Wdhx84);
	assign Kk7x84 = (Eapx84 ? Tdkw84 : L5gx84);
	assign Ek7x84 = (Eapx84 ? Ofkw84 : F9gx84);
	assign Yj7x84 = (Eapx84 ? Ailw84 : Xbgx84);
	assign Sj7x84 = (Eapx84 ? Yulw84 : Q4gx84);
	assign Mj7x84 = (Eapx84 ? Uwlw84 : E5gx84);
	assign Gj7x84 = (Lapx84 ? Kwyw84 : E5gx84);
	assign Aj7x84 = (Lapx84 ? Ouyw84 : Q4gx84);
	assign Ui7x84 = (Lapx84 ? Qhyw84 : Xbgx84);
	assign Oi7x84 = (Lapx84 ? Efxw84 : F9gx84);
	assign Ii7x84 = (Sapx84 ? Mf0x84 : E5gx84);
	assign Ci7x84 = (Sapx84 ? Qd0x84 : Q4gx84);
	assign Wh7x84 = (Sapx84 ? S00x84 : Xbgx84);
	assign Qh7x84 = (Sapx84 ? Gyyw84 : F9gx84);
	assign Kh7x84 = (Zapx84 ? Ujaw84 : Wdhx84);
	assign Eh7x84 = (Zapx84 ? Plaw84 : L5gx84);
	assign Yg7x84 = (Zapx84 ? Knaw84 : F9gx84);
	assign Sg7x84 = (Zapx84 ? Wpbw84 : Xbgx84);
	assign Mg7x84 = (Zapx84 ? U2cw84 : Q4gx84);
	assign Gg7x84 = (Zapx84 ? Q4cw84 : E5gx84);
	assign Ag7x84 = (Gbpx84 ? M6cw84 : Wdhx84);
	assign Uf7x84 = (Gbpx84 ? H8cw84 : L5gx84);
	assign Of7x84 = (Gbpx84 ? Cacw84 : F9gx84);
	assign If7x84 = (Gbpx84 ? Ocdw84 : Xbgx84);
	assign Cf7x84 = (Gbpx84 ? Mpdw84 : Q4gx84);
	assign We7x84 = (Gbpx84 ? Irdw84 : E5gx84);
	assign Qe7x84 = (Nbpx84 ? Etdw84 : Wdhx84);
	assign Ke7x84 = (Nbpx84 ? Zudw84 : L5gx84);
	assign Ee7x84 = (Nbpx84 ? Uwdw84 : F9gx84);
	assign Yd7x84 = (Nbpx84 ? Gzew84 : Xbgx84);
	assign Sd7x84 = (Nbpx84 ? Ecfw84 : Q4gx84);
	assign Md7x84 = (Nbpx84 ? Aefw84 : E5gx84);
	assign Gd7x84 = (Ubpx84 ? Wffw84 : Wdhx84);
	assign Ad7x84 = (Ubpx84 ? Rhfw84 : L5gx84);
	assign Uc7x84 = (Ubpx84 ? Mjfw84 : F9gx84);
	assign Oc7x84 = (Ubpx84 ? Ylgw84 : Xbgx84);
	assign Ic7x84 = (Ubpx84 ? Wygw84 : Q4gx84);
	assign Cc7x84 = (Ubpx84 ? S0hw84 : E5gx84);
	assign Wb7x84 = (Bcpx84 ? O2hw84 : Wdhx84);
	assign Qb7x84 = (Bcpx84 ? J4hw84 : L5gx84);
	assign Kb7x84 = (Bcpx84 ? E6hw84 : F9gx84);
	assign Eb7x84 = (Bcpx84 ? Q8iw84 : Xbgx84);
	assign Ya7x84 = (Bcpx84 ? Oliw84 : Q4gx84);
	assign Sa7x84 = (Bcpx84 ? Kniw84 : E5gx84);
	assign Ma7x84 = (Icpx84 ? Gpiw84 : Wdhx84);
	assign Wdhx84 = (~(Pcpx84 & Wcpx84));
	assign Wcpx84 = (Ddpx84 & Kdpx84);
	assign Ddpx84 = (~(Qp63a4[0] & Rdpx84));
	assign Pcpx84 = (A5ex84 & Ydpx84);
	assign Ga7x84 = (Icpx84 ? Briw84 : L5gx84);
	assign L5gx84 = (~(Gygx84 & Fepx84));
	assign Aa7x84 = (Icpx84 ? Wsiw84 : F9gx84);
	assign F9gx84 = (~(Mepx84 & Tepx84));
	assign Tepx84 = (Afpx84 & Hfpx84);
	assign Hfpx84 = (~(Qp63a4[2] & Rdpx84));
	assign Afpx84 = (Ofpx84 & Vfpx84);
	assign Vfpx84 = (~(Cgpx84 & Lwax84));
	assign Cgpx84 = (Jgpx84 & Tf63a4);
	assign Ofpx84 = (Kdpx84 | Qgpx84);
	assign Qgpx84 = (!Yk5w84);
	assign Mepx84 = (Xgpx84 & G9kx84);
	assign Xgpx84 = (Ehpx84 & Lhpx84);
	assign Lhpx84 = (Shpx84 | Zhpx84);
	assign U97x84 = (Icpx84 ? Ivjw84 : Xbgx84);
	assign O97x84 = (Icpx84 ? G8kw84 : Q4gx84);
	assign I97x84 = (Icpx84 ? Cakw84 : E5gx84);
	assign C97x84 = (Lapx84 ? Pkxw84 : Gipx84);
	assign W87x84 = (Sapx84 ? R3zw84 : Gipx84);
	assign Q87x84 = (Zapx84 ? Vsaw84 : Gipx84);
	assign K87x84 = (Gbpx84 ? Nfcw84 : Gipx84);
	assign E87x84 = (Eapx84 ? Zkkw84 : Gipx84);
	assign Y77x84 = (X9px84 ? R7mw84 : Gipx84);
	assign S77x84 = (Q9px84 ? Junw84 : Gipx84);
	assign M77x84 = (J9px84 ? Bhpw84 : Gipx84);
	assign G77x84 = (Nbpx84 ? F2ew84 : Gipx84);
	assign A77x84 = (Ubpx84 ? Xofw84 : Gipx84);
	assign U67x84 = (Bcpx84 ? Pbhw84 : Gipx84);
	assign O67x84 = (Icpx84 ? Hyiw84 : Gipx84);
	assign I67x84 = (C9px84 ? T3rw84 : Gipx84);
	assign C67x84 = (Gjhx84 ? Lqsw84 : Gipx84);
	assign W57x84 = (V8px84 ? Dduw84 : Gipx84);
	assign Q57x84 = (X4gx84 ? Vzvw84 : Gipx84);
	assign Gipx84 = (~(U2kx84 & Nipx84));
	assign K57x84 = (~(Uipx84 & Bjpx84));
	assign Bjpx84 = (Ijpx84 & Pjpx84);
	assign Pjpx84 = (~(Czdx84 & Nj63a4[5]));
	assign Ijpx84 = (~(Jzdx84 & HADDR[5]));
	assign Uipx84 = (Wjpx84 & Dkpx84);
	assign Dkpx84 = (~(Tk63a4[4] & E0ex84));
	assign Wjpx84 = (~(D69w84 & L0ex84));
	assign E57x84 = (Lapx84 ? Zgxw84 : Kkpx84);
	assign Y47x84 = (Sapx84 ? B0zw84 : Kkpx84);
	assign S47x84 = (Zapx84 ? Fpaw84 : Kkpx84);
	assign M47x84 = (Gbpx84 ? Xbcw84 : Kkpx84);
	assign G47x84 = (Eapx84 ? Jhkw84 : Kkpx84);
	assign A47x84 = (X9px84 ? B4mw84 : Kkpx84);
	assign U37x84 = (Q9px84 ? Tqnw84 : Kkpx84);
	assign O37x84 = (J9px84 ? Ldpw84 : Kkpx84);
	assign I37x84 = (Nbpx84 ? Pydw84 : Kkpx84);
	assign C37x84 = (Ubpx84 ? Hlfw84 : Kkpx84);
	assign W27x84 = (Bcpx84 ? Z7hw84 : Kkpx84);
	assign Q27x84 = (Icpx84 ? Ruiw84 : Kkpx84);
	assign K27x84 = (C9px84 ? D0rw84 : Kkpx84);
	assign E27x84 = (Gjhx84 ? Vmsw84 : Kkpx84);
	assign Y17x84 = (V8px84 ? N9uw84 : Kkpx84);
	assign S17x84 = (X4gx84 ? Fwvw84 : Kkpx84);
	assign Kkpx84 = (~(Rkpx84 & Ykpx84));
	assign Ykpx84 = (Flpx84 & Mlpx84);
	assign Mlpx84 = (Shpx84 | Tlpx84);
	assign Flpx84 = (Ampx84 & Hmpx84);
	assign Hmpx84 = (Kdpx84 | W7gx84);
	assign Ampx84 = (~(Qp63a4[3] & Rdpx84));
	assign Rkpx84 = (Tmhx84 & Ompx84);
	assign M17x84 = (~(Vmpx84 & Cnpx84));
	assign Cnpx84 = (Jnpx84 & Qnpx84);
	assign Qnpx84 = (~(Czdx84 & Nj63a4[3]));
	assign Jnpx84 = (~(Jzdx84 & HADDR[3]));
	assign Vmpx84 = (Xnpx84 & Eopx84);
	assign Eopx84 = (~(E0ex84 & Tk63a4[2]));
	assign Xnpx84 = (~(N29w84 & L0ex84));
	assign G17x84 = (~(Lopx84 & Sopx84));
	assign Sopx84 = (Zopx84 & Gppx84);
	assign Gppx84 = (~(Cr63a4[10] & Hrdx84));
	assign Zopx84 = (Nppx84 & Uppx84);
	assign Uppx84 = (Igex84 | Bqpx84);
	assign Nppx84 = (~(Qp63a4[11] & Kpdx84));
	assign Lopx84 = (Wgex84 & Iqpx84);
	assign Iqpx84 = (~(Tk63a4[10] & Ordx84));
	assign A17x84 = (~(Pqpx84 & Wqpx84));
	assign Wqpx84 = (Drpx84 & Krpx84);
	assign Krpx84 = (~(Cr63a4[18] & Hrdx84));
	assign Drpx84 = (Rrpx84 & Yrpx84);
	assign Yrpx84 = (Igex84 | Fspx84);
	assign Rrpx84 = (~(Kpdx84 & Qp63a4[19]));
	assign Pqpx84 = (Jbgx84 & Mspx84);
	assign Mspx84 = (~(Tk63a4[18] & Ordx84));
	assign U07x84 = (~(Tspx84 & Atpx84));
	assign Atpx84 = (Htpx84 & Otpx84);
	assign Otpx84 = (~(Qp63a4[27] & Kpdx84));
	assign Htpx84 = (Vtpx84 & Ypdx84);
	assign Vtpx84 = (Igex84 | Cupx84);
	assign Tspx84 = (Jupx84 & Qupx84);
	assign Qupx84 = (~(Cr63a4[26] & Hrdx84));
	assign Jupx84 = (~(Tk63a4[26] & Ordx84));
	assign O07x84 = (~(Xupx84 & Evpx84));
	assign Evpx84 = (Lvpx84 & Svpx84);
	assign Svpx84 = (~(Kpdx84 & Qp63a4[6]));
	assign Lvpx84 = (Zvpx84 & Ypdx84);
	assign Zvpx84 = (Igex84 | Gwpx84);
	assign Xupx84 = (Nwpx84 & Uwpx84);
	assign Uwpx84 = (~(Cr63a4[5] & Hrdx84));
	assign Nwpx84 = (~(Tk63a4[5] & Ordx84));
	assign I07x84 = (Lapx84 ? Kmxw84 : Bxpx84);
	assign C07x84 = (Sapx84 ? M5zw84 : Bxpx84);
	assign Wz6x84 = (Zapx84 ? Quaw84 : Bxpx84);
	assign Qz6x84 = (Gbpx84 ? Ihcw84 : Bxpx84);
	assign Kz6x84 = (Eapx84 ? Umkw84 : Bxpx84);
	assign Ez6x84 = (X9px84 ? M9mw84 : Bxpx84);
	assign Yy6x84 = (Q9px84 ? Ewnw84 : Bxpx84);
	assign Sy6x84 = (J9px84 ? Wipw84 : Bxpx84);
	assign My6x84 = (Nbpx84 ? A4ew84 : Bxpx84);
	assign Gy6x84 = (Ubpx84 ? Sqfw84 : Bxpx84);
	assign Ay6x84 = (Bcpx84 ? Kdhw84 : Bxpx84);
	assign Ux6x84 = (Icpx84 ? C0jw84 : Bxpx84);
	assign Ox6x84 = (C9px84 ? O5rw84 : Bxpx84);
	assign Ix6x84 = (Gjhx84 ? Gssw84 : Bxpx84);
	assign Cx6x84 = (V8px84 ? Yeuw84 : Bxpx84);
	assign Ww6x84 = (X4gx84 ? Q1ww84 : Bxpx84);
	assign Bxpx84 = (~(Gwpx84 & Ixpx84));
	assign Gwpx84 = (Pxpx84 & Wxpx84);
	assign Wxpx84 = (Dypx84 & Kypx84);
	assign Kypx84 = (Rypx84 | Yypx84);
	assign Dypx84 = (Fzpx84 & Mzpx84);
	assign Mzpx84 = (Tzpx84 | A0qx84);
	assign Fzpx84 = (H0qx84 | O0qx84);
	assign Pxpx84 = (V0qx84 & C1qx84);
	assign C1qx84 = (J1qx84 | Q1qx84);
	assign Qw6x84 = (~(X1qx84 & E2qx84));
	assign E2qx84 = (L2qx84 & S2qx84);
	assign S2qx84 = (~(Cr63a4[13] & Hrdx84));
	assign L2qx84 = (Z2qx84 & G3qx84);
	assign G3qx84 = (Igex84 | N3qx84);
	assign Z2qx84 = (~(Qp63a4[14] & Kpdx84));
	assign X1qx84 = (Wgex84 & U3qx84);
	assign U3qx84 = (~(Tk63a4[13] & Ordx84));
	assign Kw6x84 = (~(B4qx84 & I4qx84));
	assign I4qx84 = (P4qx84 & W4qx84);
	assign W4qx84 = (~(Cr63a4[21] & Hrdx84));
	assign P4qx84 = (D5qx84 & K5qx84);
	assign K5qx84 = (Igex84 | R5qx84);
	assign D5qx84 = (~(Qp63a4[22] & Kpdx84));
	assign B4qx84 = (Jbgx84 & Y5qx84);
	assign Y5qx84 = (~(Tk63a4[21] & Ordx84));
	assign Ew6x84 = (~(F6qx84 & M6qx84));
	assign M6qx84 = (T6qx84 & A7qx84);
	assign A7qx84 = (~(Kpdx84 & Qp63a4[4]));
	assign T6qx84 = (H7qx84 & Ypdx84);
	assign H7qx84 = (Igex84 | O7qx84);
	assign F6qx84 = (V7qx84 & C8qx84);
	assign C8qx84 = (~(Cr63a4[3] & Hrdx84));
	assign V7qx84 = (~(Tk63a4[3] & Ordx84));
	assign Yv6x84 = (~(J8qx84 & Q8qx84));
	assign Q8qx84 = (X8qx84 & E9qx84);
	assign E9qx84 = (~(Czdx84 & Nj63a4[4]));
	assign X8qx84 = (~(Jzdx84 & HADDR[4]));
	assign J8qx84 = (L9qx84 & S9qx84);
	assign S9qx84 = (~(Tk63a4[3] & E0ex84));
	assign L9qx84 = (~(I49w84 & L0ex84));
	assign Sv6x84 = (Lapx84 ? Uixw84 : Z9qx84);
	assign Mv6x84 = (Sapx84 ? W1zw84 : Z9qx84);
	assign Gv6x84 = (Zapx84 ? Araw84 : Z9qx84);
	assign Av6x84 = (Gbpx84 ? Sdcw84 : Z9qx84);
	assign Uu6x84 = (Eapx84 ? Ejkw84 : Z9qx84);
	assign Ou6x84 = (X9px84 ? W5mw84 : Z9qx84);
	assign Iu6x84 = (Q9px84 ? Osnw84 : Z9qx84);
	assign Cu6x84 = (J9px84 ? Gfpw84 : Z9qx84);
	assign Wt6x84 = (Nbpx84 ? K0ew84 : Z9qx84);
	assign Qt6x84 = (Ubpx84 ? Cnfw84 : Z9qx84);
	assign Kt6x84 = (Bcpx84 ? U9hw84 : Z9qx84);
	assign Et6x84 = (Icpx84 ? Mwiw84 : Z9qx84);
	assign Ys6x84 = (C9px84 ? Y1rw84 : Z9qx84);
	assign Ss6x84 = (Gjhx84 ? Qosw84 : Z9qx84);
	assign Ms6x84 = (V8px84 ? Ibuw84 : Z9qx84);
	assign Gs6x84 = (X4gx84 ? Ayvw84 : Z9qx84);
	assign Z9qx84 = (~(O7qx84 & Gaqx84));
	assign As6x84 = (~(Naqx84 & Uaqx84));
	assign Uaqx84 = (Bbqx84 & Ibqx84);
	assign Ibqx84 = (~(Cr63a4[11] & Hrdx84));
	assign Bbqx84 = (Pbqx84 & Wbqx84);
	assign Wbqx84 = (Igex84 | Dcqx84);
	assign Pbqx84 = (~(Kpdx84 & Qp63a4[12]));
	assign Naqx84 = (Wgex84 & Kcqx84);
	assign Kcqx84 = (~(Tk63a4[11] & Ordx84));
	assign Wgex84 = (Rcqx84 & Ypdx84);
	assign Rcqx84 = (Ycqx84 | Igex84);
	assign Ur6x84 = (~(Fdqx84 & Mdqx84));
	assign Mdqx84 = (Tdqx84 & Aeqx84);
	assign Aeqx84 = (~(Cr63a4[19] & Hrdx84));
	assign Tdqx84 = (Heqx84 & Oeqx84);
	assign Oeqx84 = (Igex84 | Veqx84);
	assign Heqx84 = (~(Qp63a4[20] & Kpdx84));
	assign Fdqx84 = (Jbgx84 & Cfqx84);
	assign Cfqx84 = (~(Tk63a4[19] & Ordx84));
	assign Or6x84 = (~(Jfqx84 & Qfqx84));
	assign Qfqx84 = (Xfqx84 & Egqx84);
	assign Egqx84 = (~(Qp63a4[28] & Kpdx84));
	assign Xfqx84 = (Lgqx84 & Ypdx84);
	assign Lgqx84 = (Igex84 | Sgqx84);
	assign Jfqx84 = (Zgqx84 & Ghqx84);
	assign Ghqx84 = (~(Cr63a4[27] & Hrdx84));
	assign Zgqx84 = (~(Tk63a4[27] & Ordx84));
	assign Ir6x84 = (Lapx84 ? Foxw84 : Njhx84);
	assign Cr6x84 = (Sapx84 ? H7zw84 : Njhx84);
	assign Wq6x84 = (Zapx84 ? Lwaw84 : Njhx84);
	assign Qq6x84 = (Gbpx84 ? Djcw84 : Njhx84);
	assign Kq6x84 = (Eapx84 ? Pokw84 : Njhx84);
	assign Eq6x84 = (X9px84 ? Hbmw84 : Njhx84);
	assign Yp6x84 = (Q9px84 ? Zxnw84 : Njhx84);
	assign Sp6x84 = (J9px84 ? Rkpw84 : Njhx84);
	assign Mp6x84 = (Nbpx84 ? V5ew84 : Njhx84);
	assign Gp6x84 = (Ubpx84 ? Nsfw84 : Njhx84);
	assign Ap6x84 = (Bcpx84 ? Ffhw84 : Njhx84);
	assign Uo6x84 = (Icpx84 ? X1jw84 : Njhx84);
	assign Oo6x84 = (C9px84 ? J7rw84 : Njhx84);
	assign Io6x84 = (V8px84 ? Tguw84 : Njhx84);
	assign Co6x84 = (X4gx84 ? L3ww84 : Njhx84);
	assign Njhx84 = (~(Nhqx84 & Uhqx84));
	assign Uhqx84 = (Biqx84 & Iiqx84);
	assign Iiqx84 = (Shpx84 | Piqx84);
	assign Biqx84 = (Wiqx84 & Kdpx84);
	assign Wiqx84 = (~(Qp63a4[7] & Rdpx84));
	assign Nhqx84 = (~(Djqx84 | Kyix84));
	assign Kyix84 = (~(Kjqx84 & Rjqx84));
	assign Rjqx84 = (Yjqx84 & Fkqx84);
	assign Fkqx84 = (J1qx84 | Mkqx84);
	assign Yjqx84 = (Tkqx84 & Alqx84);
	assign Alqx84 = (H0qx84 | Hlqx84);
	assign Tkqx84 = (Rypx84 | Olqx84);
	assign Kjqx84 = (V0qx84 & Vlqx84);
	assign Vlqx84 = (Tzpx84 | Cmqx84);
	assign Djqx84 = (Ftax84 ? Qmqx84 : Jmqx84);
	assign Qmqx84 = (Jgpx84 & Gj63a4);
	assign Wn6x84 = (Gjhx84 ? Wvsw84 : Xmqx84);
	assign Qn6x84 = (Lapx84 ? Aqxw84 : Xmqx84);
	assign Kn6x84 = (Sapx84 ? C9zw84 : Xmqx84);
	assign En6x84 = (Zapx84 ? Gyaw84 : Xmqx84);
	assign Ym6x84 = (Gbpx84 ? Ykcw84 : Xmqx84);
	assign Sm6x84 = (Eapx84 ? Kqkw84 : Xmqx84);
	assign Mm6x84 = (X9px84 ? Cdmw84 : Xmqx84);
	assign Gm6x84 = (Q9px84 ? Uznw84 : Xmqx84);
	assign Am6x84 = (J9px84 ? Mmpw84 : Xmqx84);
	assign Ul6x84 = (Nbpx84 ? Q7ew84 : Xmqx84);
	assign Ol6x84 = (Ubpx84 ? Iufw84 : Xmqx84);
	assign Il6x84 = (Bcpx84 ? Ahhw84 : Xmqx84);
	assign Cl6x84 = (Icpx84 ? S3jw84 : Xmqx84);
	assign Wk6x84 = (C9px84 ? E9rw84 : Xmqx84);
	assign Qk6x84 = (V8px84 ? Oiuw84 : Xmqx84);
	assign Kk6x84 = (X4gx84 ? G5ww84 : Xmqx84);
	assign Xmqx84 = (~(Enqx84 & Pgex84));
	assign Pgex84 = (Lnqx84 & Snqx84);
	assign Snqx84 = (Znqx84 & Goqx84);
	assign Goqx84 = (Noqx84 | Uoqx84);
	assign Znqx84 = (Bpqx84 | Ipqx84);
	assign Lnqx84 = (Ppqx84 & Wpqx84);
	assign Wpqx84 = (Dqqx84 | Kqqx84);
	assign Ppqx84 = (Rqqx84 | Yqqx84);
	assign Enqx84 = (Frqx84 & Ycqx84);
	assign Ek6x84 = (Gjhx84 ? Rxsw84 : Mrqx84);
	assign Yj6x84 = (Lapx84 ? Vrxw84 : Mrqx84);
	assign Sj6x84 = (Sapx84 ? Xazw84 : Mrqx84);
	assign Mj6x84 = (Zapx84 ? B0bw84 : Mrqx84);
	assign Gj6x84 = (Gbpx84 ? Tmcw84 : Mrqx84);
	assign Aj6x84 = (Eapx84 ? Fskw84 : Mrqx84);
	assign Ui6x84 = (X9px84 ? Xemw84 : Mrqx84);
	assign Oi6x84 = (Q9px84 ? P1ow84 : Mrqx84);
	assign Ii6x84 = (J9px84 ? Hopw84 : Mrqx84);
	assign Ci6x84 = (Nbpx84 ? L9ew84 : Mrqx84);
	assign Wh6x84 = (Ubpx84 ? Dwfw84 : Mrqx84);
	assign Qh6x84 = (Bcpx84 ? Vihw84 : Mrqx84);
	assign Kh6x84 = (Icpx84 ? N5jw84 : Mrqx84);
	assign Eh6x84 = (C9px84 ? Zarw84 : Mrqx84);
	assign Yg6x84 = (V8px84 ? Jkuw84 : Mrqx84);
	assign Sg6x84 = (X4gx84 ? B7ww84 : Mrqx84);
	assign Mrqx84 = (~(Bpcx84 & Trqx84));
	assign Bpcx84 = (Asqx84 & Hsqx84);
	assign Hsqx84 = (Osqx84 & Vsqx84);
	assign Vsqx84 = (Ipqx84 | Ctqx84);
	assign Osqx84 = (Jtqx84 & Ycqx84);
	assign Jtqx84 = (Uoqx84 | Qtqx84);
	assign Asqx84 = (Xtqx84 & Euqx84);
	assign Euqx84 = (Kqqx84 | Luqx84);
	assign Xtqx84 = (Yqqx84 | Suqx84);
	assign Mg6x84 = (Gjhx84 ? Mzsw84 : Zuqx84);
	assign Gg6x84 = (Lapx84 ? Qtxw84 : Zuqx84);
	assign Ag6x84 = (Sapx84 ? Sczw84 : Zuqx84);
	assign Uf6x84 = (Zapx84 ? W1bw84 : Zuqx84);
	assign Of6x84 = (Gbpx84 ? Oocw84 : Zuqx84);
	assign If6x84 = (Eapx84 ? Aukw84 : Zuqx84);
	assign Cf6x84 = (X9px84 ? Sgmw84 : Zuqx84);
	assign We6x84 = (Q9px84 ? K3ow84 : Zuqx84);
	assign Qe6x84 = (J9px84 ? Cqpw84 : Zuqx84);
	assign Ke6x84 = (Nbpx84 ? Gbew84 : Zuqx84);
	assign Ee6x84 = (Ubpx84 ? Yxfw84 : Zuqx84);
	assign Yd6x84 = (Bcpx84 ? Qkhw84 : Zuqx84);
	assign Sd6x84 = (Icpx84 ? I7jw84 : Zuqx84);
	assign Md6x84 = (C9px84 ? Ucrw84 : Zuqx84);
	assign Gd6x84 = (V8px84 ? Emuw84 : Zuqx84);
	assign Ad6x84 = (X4gx84 ? W8ww84 : Zuqx84);
	assign Zuqx84 = (~(Gvqx84 & Nvqx84));
	assign Nvqx84 = (Uvqx84 & Bwqx84);
	assign Bwqx84 = (~(Qp63a4[10] & Rdpx84));
	assign Uvqx84 = (Iwqx84 & Pwqx84);
	assign Iwqx84 = (~(Wwqx84 & C2bx84));
	assign Wwqx84 = (Jgpx84 & Xh63a4);
	assign Gvqx84 = (Dxqx84 & Kxqx84);
	assign Dxqx84 = (Rbkx84 & Rxqx84);
	assign Rxqx84 = (Shpx84 | Yxqx84);
	assign Rbkx84 = (Fyqx84 & Myqx84);
	assign Myqx84 = (Tyqx84 & Azqx84);
	assign Azqx84 = (Hzqx84 | Uoqx84);
	assign Tyqx84 = (Ozqx84 | Ipqx84);
	assign Fyqx84 = (Vzqx84 & C0rx84);
	assign C0rx84 = (J0rx84 | Kqqx84);
	assign Vzqx84 = (Q0rx84 | Yqqx84);
	assign Uc6x84 = (Gjhx84 ? I1tw84 : X0rx84);
	assign Oc6x84 = (Lapx84 ? Mvxw84 : X0rx84);
	assign Ic6x84 = (Sapx84 ? Oezw84 : X0rx84);
	assign Cc6x84 = (Zapx84 ? S3bw84 : X0rx84);
	assign Wb6x84 = (Gbpx84 ? Kqcw84 : X0rx84);
	assign Qb6x84 = (Eapx84 ? Wvkw84 : X0rx84);
	assign Kb6x84 = (X9px84 ? Oimw84 : X0rx84);
	assign Eb6x84 = (Q9px84 ? G5ow84 : X0rx84);
	assign Ya6x84 = (J9px84 ? Yrpw84 : X0rx84);
	assign Sa6x84 = (Nbpx84 ? Cdew84 : X0rx84);
	assign Ma6x84 = (Ubpx84 ? Uzfw84 : X0rx84);
	assign Ga6x84 = (Bcpx84 ? Mmhw84 : X0rx84);
	assign Aa6x84 = (Icpx84 ? E9jw84 : X0rx84);
	assign U96x84 = (C9px84 ? Qerw84 : X0rx84);
	assign O96x84 = (V8px84 ? Aouw84 : X0rx84);
	assign I96x84 = (X4gx84 ? Saww84 : X0rx84);
	assign X0rx84 = (~(E1rx84 & L1rx84));
	assign L1rx84 = (S1rx84 & Z1rx84);
	assign Z1rx84 = (~(Qp63a4[11] & Rdpx84));
	assign S1rx84 = (G2rx84 & N2rx84);
	assign G2rx84 = (~(U2rx84 & V1bx84));
	assign U2rx84 = (Jgpx84 & Zi63a4);
	assign E1rx84 = (B3rx84 & Bqpx84);
	assign Bqpx84 = (I3rx84 & P3rx84);
	assign P3rx84 = (W3rx84 & D4rx84);
	assign D4rx84 = (K4rx84 | Uoqx84);
	assign W3rx84 = (R4rx84 | Ipqx84);
	assign I3rx84 = (Y4rx84 & F5rx84);
	assign F5rx84 = (M5rx84 | Kqqx84);
	assign Y4rx84 = (T5rx84 | Yqqx84);
	assign B3rx84 = (Kxqx84 & A6rx84);
	assign A6rx84 = (Shpx84 | H6rx84);
	assign C96x84 = (Gjhx84 ? E3tw84 : O6rx84);
	assign W86x84 = (Lapx84 ? Ixxw84 : O6rx84);
	assign Q86x84 = (Sapx84 ? Kgzw84 : O6rx84);
	assign K86x84 = (Zapx84 ? O5bw84 : O6rx84);
	assign E86x84 = (Gbpx84 ? Gscw84 : O6rx84);
	assign Y76x84 = (Eapx84 ? Sxkw84 : O6rx84);
	assign S76x84 = (X9px84 ? Kkmw84 : O6rx84);
	assign M76x84 = (Q9px84 ? C7ow84 : O6rx84);
	assign G76x84 = (J9px84 ? Utpw84 : O6rx84);
	assign A76x84 = (Nbpx84 ? Yeew84 : O6rx84);
	assign U66x84 = (Ubpx84 ? Q1gw84 : O6rx84);
	assign O66x84 = (Bcpx84 ? Iohw84 : O6rx84);
	assign I66x84 = (Icpx84 ? Abjw84 : O6rx84);
	assign C66x84 = (C9px84 ? Mgrw84 : O6rx84);
	assign W56x84 = (V8px84 ? Wpuw84 : O6rx84);
	assign Q56x84 = (X4gx84 ? Ocww84 : O6rx84);
	assign O6rx84 = (~(V6rx84 & Dcqx84));
	assign Dcqx84 = (C7rx84 & J7rx84);
	assign J7rx84 = (Q7rx84 & X7rx84);
	assign X7rx84 = (E8rx84 | Uoqx84);
	assign Q7rx84 = (L8rx84 | Ipqx84);
	assign C7rx84 = (S8rx84 & Z8rx84);
	assign Z8rx84 = (G9rx84 | Kqqx84);
	assign S8rx84 = (N9rx84 | Yqqx84);
	assign V6rx84 = (U9rx84 & Ycqx84);
	assign K56x84 = (Gjhx84 ? A5tw84 : Barx84);
	assign E56x84 = (Lapx84 ? Ezxw84 : Barx84);
	assign Y46x84 = (Sapx84 ? Gizw84 : Barx84);
	assign S46x84 = (Zapx84 ? K7bw84 : Barx84);
	assign M46x84 = (Gbpx84 ? Cucw84 : Barx84);
	assign G46x84 = (Eapx84 ? Ozkw84 : Barx84);
	assign A46x84 = (X9px84 ? Gmmw84 : Barx84);
	assign U36x84 = (Q9px84 ? Y8ow84 : Barx84);
	assign O36x84 = (J9px84 ? Qvpw84 : Barx84);
	assign I36x84 = (Nbpx84 ? Ugew84 : Barx84);
	assign C36x84 = (Ubpx84 ? M3gw84 : Barx84);
	assign W26x84 = (Bcpx84 ? Eqhw84 : Barx84);
	assign Q26x84 = (Icpx84 ? Wcjw84 : Barx84);
	assign K26x84 = (C9px84 ? Iirw84 : Barx84);
	assign E26x84 = (V8px84 ? Sruw84 : Barx84);
	assign Y16x84 = (X4gx84 ? Keww84 : Barx84);
	assign Barx84 = (~(Iarx84 & Parx84));
	assign Parx84 = (Warx84 & Dbrx84);
	assign Dbrx84 = (~(Qp63a4[13] & Rdpx84));
	assign Warx84 = (Kbrx84 & Rbrx84);
	assign Kbrx84 = (~(Ybrx84 & H1bx84));
	assign Ybrx84 = (Jgpx84 & Ei63a4);
	assign Iarx84 = (Fcrx84 & F5kx84);
	assign F5kx84 = (Mcrx84 & Tcrx84);
	assign Tcrx84 = (Adrx84 & Hdrx84);
	assign Hdrx84 = (Odrx84 | Uoqx84);
	assign Adrx84 = (Vdrx84 | Ipqx84);
	assign Mcrx84 = (Cerx84 & Jerx84);
	assign Jerx84 = (Qerx84 | Kqqx84);
	assign Cerx84 = (Xerx84 | Yqqx84);
	assign Fcrx84 = (Kxqx84 & Efrx84);
	assign Efrx84 = (Shpx84 | Lfrx84);
	assign S16x84 = (Gjhx84 ? W6tw84 : Sfrx84);
	assign M16x84 = (Lapx84 ? A1yw84 : Sfrx84);
	assign G16x84 = (Sapx84 ? Ckzw84 : Sfrx84);
	assign A16x84 = (Zapx84 ? G9bw84 : Sfrx84);
	assign U06x84 = (Gbpx84 ? Yvcw84 : Sfrx84);
	assign O06x84 = (Eapx84 ? K1lw84 : Sfrx84);
	assign I06x84 = (X9px84 ? Comw84 : Sfrx84);
	assign C06x84 = (Q9px84 ? Uaow84 : Sfrx84);
	assign Wz5x84 = (J9px84 ? Mxpw84 : Sfrx84);
	assign Qz5x84 = (Nbpx84 ? Qiew84 : Sfrx84);
	assign Kz5x84 = (Ubpx84 ? I5gw84 : Sfrx84);
	assign Ez5x84 = (Bcpx84 ? Ashw84 : Sfrx84);
	assign Yy5x84 = (Icpx84 ? Sejw84 : Sfrx84);
	assign Sy5x84 = (C9px84 ? Ekrw84 : Sfrx84);
	assign My5x84 = (V8px84 ? Otuw84 : Sfrx84);
	assign Gy5x84 = (X4gx84 ? Ggww84 : Sfrx84);
	assign Sfrx84 = (~(Zfrx84 & Ggrx84));
	assign Ggrx84 = (Ngrx84 & Ugrx84);
	assign Ugrx84 = (~(Qp63a4[14] & Rdpx84));
	assign Ngrx84 = (Bhrx84 & Ihrx84);
	assign Bhrx84 = (~(Phrx84 & A1bx84));
	assign Phrx84 = (Jgpx84 & Li63a4);
	assign Zfrx84 = (Whrx84 & N3qx84);
	assign N3qx84 = (Dirx84 & Kirx84);
	assign Kirx84 = (Rirx84 & Yirx84);
	assign Yirx84 = (Q1qx84 | Uoqx84);
	assign Rirx84 = (Yypx84 | Ipqx84);
	assign Dirx84 = (Fjrx84 & Mjrx84);
	assign Mjrx84 = (O0qx84 | Kqqx84);
	assign Fjrx84 = (A0qx84 | Yqqx84);
	assign Whrx84 = (Kxqx84 & Tjrx84);
	assign Tjrx84 = (Shpx84 | Akrx84);
	assign Ay5x84 = (Gjhx84 ? S8tw84 : Hkrx84);
	assign Ux5x84 = (Lapx84 ? W2yw84 : Hkrx84);
	assign Ox5x84 = (Sapx84 ? Ylzw84 : Hkrx84);
	assign Ix5x84 = (Zapx84 ? Cbbw84 : Hkrx84);
	assign Cx5x84 = (Gbpx84 ? Uxcw84 : Hkrx84);
	assign Ww5x84 = (Eapx84 ? G3lw84 : Hkrx84);
	assign Qw5x84 = (X9px84 ? Ypmw84 : Hkrx84);
	assign Kw5x84 = (Q9px84 ? Qcow84 : Hkrx84);
	assign Ew5x84 = (J9px84 ? Izpw84 : Hkrx84);
	assign Yv5x84 = (Nbpx84 ? Mkew84 : Hkrx84);
	assign Sv5x84 = (Ubpx84 ? E7gw84 : Hkrx84);
	assign Mv5x84 = (Bcpx84 ? Wthw84 : Hkrx84);
	assign Gv5x84 = (Icpx84 ? Ogjw84 : Hkrx84);
	assign Av5x84 = (C9px84 ? Amrw84 : Hkrx84);
	assign Uu5x84 = (V8px84 ? Kvuw84 : Hkrx84);
	assign Ou5x84 = (X4gx84 ? Ciww84 : Hkrx84);
	assign Hkrx84 = (~(Okrx84 & Vkrx84));
	assign Vkrx84 = (Clrx84 & Jlrx84);
	assign Jlrx84 = (~(Qp63a4[15] & Rdpx84));
	assign Clrx84 = (Qlrx84 & Xlrx84);
	assign Qlrx84 = (~(Emrx84 & T0bx84));
	assign Emrx84 = (Jgpx84 & Si63a4);
	assign Okrx84 = (Lmrx84 & V0jx84);
	assign V0jx84 = (Smrx84 & Zmrx84);
	assign Zmrx84 = (Gnrx84 & Nnrx84);
	assign Nnrx84 = (Uoqx84 | Mkqx84);
	assign Uoqx84 = (Unrx84 & Borx84);
	assign Gnrx84 = (Ipqx84 | Olqx84);
	assign Ipqx84 = (Iorx84 & Porx84);
	assign Porx84 = (~(Worx84 & Dprx84));
	assign Dprx84 = (Kprx84 | Ozcx84);
	assign Worx84 = (~(Rprx84 | Vs63a4[1]));
	assign Smrx84 = (Yprx84 & Fqrx84);
	assign Fqrx84 = (Kqqx84 | Hlqx84);
	assign Kqqx84 = (Mqrx84 & Tqrx84);
	assign Tqrx84 = (~(Arrx84 & Vs63a4[1]));
	assign Arrx84 = (Hrrx84 & Orrx84);
	assign Hrrx84 = (~(Bdox84 & Vrrx84));
	assign Vrrx84 = (~(Csrx84 & Jsrx84));
	assign Csrx84 = (~(Hu2x84 | J13x84));
	assign Yprx84 = (Yqqx84 | Cmqx84);
	assign Yqqx84 = (Qsrx84 & Xsrx84);
	assign Lmrx84 = (Kxqx84 & Etrx84);
	assign Etrx84 = (Shpx84 | Ltrx84);
	assign Kxqx84 = (Kdpx84 & Ycqx84);
	assign Ycqx84 = (~(Strx84 & Ztrx84));
	assign Ztrx84 = (Gurx84 & Xsrx84);
	assign Strx84 = (Nurx84 & Mqrx84);
	assign Nurx84 = (Orrx84 ? Bvrx84 : Uurx84);
	assign Bvrx84 = (~(Ivrx84 & Pvrx84));
	assign Iu5x84 = (Gjhx84 ? Kctw84 : Wvrx84);
	assign Cu5x84 = (Lapx84 ? O6yw84 : Wvrx84);
	assign Wt5x84 = (Sapx84 ? Qpzw84 : Wvrx84);
	assign Qt5x84 = (Zapx84 ? Uebw84 : Wvrx84);
	assign Kt5x84 = (Gbpx84 ? M1dw84 : Wvrx84);
	assign Et5x84 = (Eapx84 ? Y6lw84 : Wvrx84);
	assign Ys5x84 = (X9px84 ? Qtmw84 : Wvrx84);
	assign Ss5x84 = (Q9px84 ? Igow84 : Wvrx84);
	assign Ms5x84 = (J9px84 ? A3qw84 : Wvrx84);
	assign Gs5x84 = (Nbpx84 ? Eoew84 : Wvrx84);
	assign As5x84 = (Ubpx84 ? Wagw84 : Wvrx84);
	assign Ur5x84 = (Bcpx84 ? Oxhw84 : Wvrx84);
	assign Or5x84 = (Icpx84 ? Gkjw84 : Wvrx84);
	assign Ir5x84 = (C9px84 ? Sprw84 : Wvrx84);
	assign Cr5x84 = (V8px84 ? Czuw84 : Wvrx84);
	assign Wq5x84 = (X4gx84 ? Ulww84 : Wvrx84);
	assign Wvrx84 = (~(Dwrx84 & Dxjx84));
	assign Dxjx84 = (Kwrx84 & Rwrx84);
	assign Rwrx84 = (Ywrx84 & Fxrx84);
	assign Fxrx84 = (Mxrx84 | Ctqx84);
	assign Ywrx84 = (Txrx84 | Luqx84);
	assign Kwrx84 = (Ayrx84 & Hyrx84);
	assign Hyrx84 = (Oyrx84 | Suqx84);
	assign Ayrx84 = (Vyrx84 | Qtqx84);
	assign Dwrx84 = (Czrx84 & Jzrx84);
	assign Qq5x84 = (Gjhx84 ? Getw84 : Qzrx84);
	assign Kq5x84 = (Lapx84 ? K8yw84 : Qzrx84);
	assign Eq5x84 = (Sapx84 ? Mrzw84 : Qzrx84);
	assign Yp5x84 = (Zapx84 ? Qgbw84 : Qzrx84);
	assign Sp5x84 = (Gbpx84 ? I3dw84 : Qzrx84);
	assign Mp5x84 = (Eapx84 ? U8lw84 : Qzrx84);
	assign Gp5x84 = (X9px84 ? Mvmw84 : Qzrx84);
	assign Ap5x84 = (Q9px84 ? Eiow84 : Qzrx84);
	assign Uo5x84 = (J9px84 ? W4qw84 : Qzrx84);
	assign Oo5x84 = (Nbpx84 ? Aqew84 : Qzrx84);
	assign Io5x84 = (Ubpx84 ? Scgw84 : Qzrx84);
	assign Co5x84 = (Bcpx84 ? Kzhw84 : Qzrx84);
	assign Wn5x84 = (Icpx84 ? Cmjw84 : Qzrx84);
	assign Qn5x84 = (C9px84 ? Orrw84 : Qzrx84);
	assign Kn5x84 = (V8px84 ? Y0vw84 : Qzrx84);
	assign En5x84 = (X4gx84 ? Qnww84 : Qzrx84);
	assign Qzrx84 = (~(Xzrx84 & Vdkx84));
	assign Vdkx84 = (E0sx84 & L0sx84);
	assign L0sx84 = (S0sx84 & Z0sx84);
	assign Z0sx84 = (Mxrx84 | Ozqx84);
	assign S0sx84 = (Txrx84 | J0rx84);
	assign E0sx84 = (G1sx84 & N1sx84);
	assign N1sx84 = (Oyrx84 | Q0rx84);
	assign G1sx84 = (Vyrx84 | Hzqx84);
	assign Xzrx84 = (Czrx84 & U1sx84);
	assign Ym5x84 = (Gjhx84 ? Cgtw84 : B2sx84);
	assign Sm5x84 = (Lapx84 ? Gayw84 : B2sx84);
	assign Mm5x84 = (Sapx84 ? Itzw84 : B2sx84);
	assign Gm5x84 = (Zapx84 ? Mibw84 : B2sx84);
	assign Am5x84 = (Gbpx84 ? E5dw84 : B2sx84);
	assign Ul5x84 = (Eapx84 ? Qalw84 : B2sx84);
	assign Ol5x84 = (X9px84 ? Ixmw84 : B2sx84);
	assign Il5x84 = (Q9px84 ? Akow84 : B2sx84);
	assign Cl5x84 = (J9px84 ? S6qw84 : B2sx84);
	assign Wk5x84 = (Nbpx84 ? Wrew84 : B2sx84);
	assign Qk5x84 = (Ubpx84 ? Oegw84 : B2sx84);
	assign Kk5x84 = (Bcpx84 ? G1iw84 : B2sx84);
	assign Ek5x84 = (Icpx84 ? Ynjw84 : B2sx84);
	assign Yj5x84 = (C9px84 ? Ktrw84 : B2sx84);
	assign Sj5x84 = (V8px84 ? U2vw84 : B2sx84);
	assign Mj5x84 = (X4gx84 ? Mpww84 : B2sx84);
	assign B2sx84 = (~(I2sx84 & Fspx84));
	assign Fspx84 = (P2sx84 & W2sx84);
	assign W2sx84 = (D3sx84 & K3sx84);
	assign K3sx84 = (R4rx84 | Mxrx84);
	assign D3sx84 = (Txrx84 | M5rx84);
	assign P2sx84 = (R3sx84 & Y3sx84);
	assign Y3sx84 = (Oyrx84 | T5rx84);
	assign R3sx84 = (Vyrx84 | K4rx84);
	assign I2sx84 = (Czrx84 & F4sx84);
	assign Gj5x84 = (Gjhx84 ? Yhtw84 : M4sx84);
	assign Aj5x84 = (Lapx84 ? Ccyw84 : M4sx84);
	assign Ui5x84 = (Sapx84 ? Evzw84 : M4sx84);
	assign Oi5x84 = (Zapx84 ? Ikbw84 : M4sx84);
	assign Ii5x84 = (Gbpx84 ? A7dw84 : M4sx84);
	assign Ci5x84 = (Eapx84 ? Mclw84 : M4sx84);
	assign Wh5x84 = (X9px84 ? Ezmw84 : M4sx84);
	assign Qh5x84 = (Q9px84 ? Wlow84 : M4sx84);
	assign Kh5x84 = (J9px84 ? O8qw84 : M4sx84);
	assign Eh5x84 = (Nbpx84 ? Stew84 : M4sx84);
	assign Yg5x84 = (Ubpx84 ? Kggw84 : M4sx84);
	assign Sg5x84 = (Bcpx84 ? C3iw84 : M4sx84);
	assign Mg5x84 = (Icpx84 ? Upjw84 : M4sx84);
	assign Gg5x84 = (C9px84 ? Gvrw84 : M4sx84);
	assign Ag5x84 = (V8px84 ? Q4vw84 : M4sx84);
	assign Uf5x84 = (X4gx84 ? Irww84 : M4sx84);
	assign M4sx84 = (~(T4sx84 & A5sx84));
	assign A5sx84 = (H5sx84 & O5sx84);
	assign O5sx84 = (~(Qp63a4[20] & Rdpx84));
	assign H5sx84 = (V5sx84 & C6sx84);
	assign V5sx84 = (~(J6sx84 & Dzax84));
	assign J6sx84 = (Jgpx84 & Og63a4);
	assign T4sx84 = (Q6sx84 & Veqx84);
	assign Veqx84 = (X6sx84 & E7sx84);
	assign E7sx84 = (L7sx84 & S7sx84);
	assign S7sx84 = (L8rx84 | Mxrx84);
	assign L7sx84 = (Txrx84 | G9rx84);
	assign X6sx84 = (Z7sx84 & G8sx84);
	assign G8sx84 = (Oyrx84 | N9rx84);
	assign Z7sx84 = (Vyrx84 | E8rx84);
	assign Q6sx84 = (N8sx84 & U8sx84);
	assign U8sx84 = (Shpx84 | B9sx84);
	assign Of5x84 = (Gjhx84 ? Ujtw84 : I9sx84);
	assign If5x84 = (Lapx84 ? Ydyw84 : I9sx84);
	assign Cf5x84 = (Sapx84 ? Axzw84 : I9sx84);
	assign We5x84 = (Zapx84 ? Embw84 : I9sx84);
	assign Qe5x84 = (Gbpx84 ? W8dw84 : I9sx84);
	assign Ke5x84 = (Eapx84 ? Ielw84 : I9sx84);
	assign Ee5x84 = (X9px84 ? A1nw84 : I9sx84);
	assign Yd5x84 = (Q9px84 ? Snow84 : I9sx84);
	assign Sd5x84 = (J9px84 ? Kaqw84 : I9sx84);
	assign Md5x84 = (Nbpx84 ? Ovew84 : I9sx84);
	assign Gd5x84 = (Ubpx84 ? Gigw84 : I9sx84);
	assign Ad5x84 = (Bcpx84 ? Y4iw84 : I9sx84);
	assign Uc5x84 = (Icpx84 ? Qrjw84 : I9sx84);
	assign Oc5x84 = (C9px84 ? Cxrw84 : I9sx84);
	assign Ic5x84 = (V8px84 ? M6vw84 : I9sx84);
	assign Cc5x84 = (X4gx84 ? Etww84 : I9sx84);
	assign I9sx84 = (~(P9sx84 & W9sx84));
	assign W9sx84 = (Dasx84 & Kasx84);
	assign Kasx84 = (~(Qp63a4[21] & Rdpx84));
	assign Dasx84 = (Rasx84 & Yasx84);
	assign Rasx84 = (~(Fbsx84 & Wyax84));
	assign Fbsx84 = (Jgpx84 & Vg63a4);
	assign P9sx84 = (Mbsx84 & J7kx84);
	assign J7kx84 = (Tbsx84 & Acsx84);
	assign Acsx84 = (Hcsx84 & Ocsx84);
	assign Ocsx84 = (Vdrx84 | Mxrx84);
	assign Hcsx84 = (Txrx84 | Qerx84);
	assign Tbsx84 = (Vcsx84 & Cdsx84);
	assign Cdsx84 = (Oyrx84 | Xerx84);
	assign Vcsx84 = (Vyrx84 | Odrx84);
	assign Mbsx84 = (N8sx84 & Jdsx84);
	assign Jdsx84 = (Shpx84 | Qdsx84);
	assign Wb5x84 = (Gjhx84 ? Qltw84 : Xdsx84);
	assign Qb5x84 = (Lapx84 ? Ufyw84 : Xdsx84);
	assign Kb5x84 = (Sapx84 ? Wyzw84 : Xdsx84);
	assign Eb5x84 = (Zapx84 ? Aobw84 : Xdsx84);
	assign Ya5x84 = (Gbpx84 ? Sadw84 : Xdsx84);
	assign Sa5x84 = (Eapx84 ? Eglw84 : Xdsx84);
	assign Ma5x84 = (X9px84 ? W2nw84 : Xdsx84);
	assign Ga5x84 = (Q9px84 ? Opow84 : Xdsx84);
	assign Aa5x84 = (J9px84 ? Gcqw84 : Xdsx84);
	assign U95x84 = (Nbpx84 ? Kxew84 : Xdsx84);
	assign O95x84 = (Ubpx84 ? Ckgw84 : Xdsx84);
	assign I95x84 = (Bcpx84 ? U6iw84 : Xdsx84);
	assign C95x84 = (Icpx84 ? Mtjw84 : Xdsx84);
	assign W85x84 = (C9px84 ? Yyrw84 : Xdsx84);
	assign Q85x84 = (V8px84 ? I8vw84 : Xdsx84);
	assign K85x84 = (X4gx84 ? Avww84 : Xdsx84);
	assign Xdsx84 = (~(Eesx84 & Lesx84));
	assign Lesx84 = (Sesx84 & Zesx84);
	assign Zesx84 = (~(Qp63a4[22] & Rdpx84));
	assign Sesx84 = (Gfsx84 & Nfsx84);
	assign Gfsx84 = (~(Ufsx84 & Pyax84));
	assign Ufsx84 = (Jgpx84 & Jh63a4);
	assign Eesx84 = (Bgsx84 & R5qx84);
	assign R5qx84 = (Igsx84 & Pgsx84);
	assign Pgsx84 = (Wgsx84 & Dhsx84);
	assign Dhsx84 = (Oyrx84 | A0qx84);
	assign Wgsx84 = (Txrx84 | O0qx84);
	assign Igsx84 = (Khsx84 & Rhsx84);
	assign Rhsx84 = (Mxrx84 | Yypx84);
	assign Khsx84 = (Vyrx84 | Q1qx84);
	assign Bgsx84 = (N8sx84 & Yhsx84);
	assign Yhsx84 = (Shpx84 | Fisx84);
	assign E85x84 = (Gjhx84 ? Mntw84 : Xbgx84);
	assign Xbgx84 = (~(Misx84 & Tisx84));
	assign Tisx84 = (Ajsx84 & Hjsx84);
	assign Hjsx84 = (~(Qp63a4[23] & Rdpx84));
	assign Ajsx84 = (Ojsx84 & Vjsx84);
	assign Ojsx84 = (~(Cksx84 & Iyax84));
	assign Cksx84 = (Jgpx84 & Qh63a4);
	assign Misx84 = (Jksx84 & N8sx84);
	assign Jksx84 = (Cbgx84 & Qksx84);
	assign Qksx84 = (Shpx84 | Xksx84);
	assign Cbgx84 = (Elsx84 & Llsx84);
	assign Llsx84 = (Slsx84 & Zlsx84);
	assign Zlsx84 = (Mxrx84 | Olqx84);
	assign Slsx84 = (Txrx84 | Hlqx84);
	assign Elsx84 = (Gmsx84 & Nmsx84);
	assign Nmsx84 = (Oyrx84 | Cmqx84);
	assign Gmsx84 = (Vyrx84 | Mkqx84);
	assign Y75x84 = (Gjhx84 ? Ertw84 : Umsx84);
	assign S75x84 = (Lapx84 ? Ilyw84 : Umsx84);
	assign M75x84 = (Sapx84 ? K40x84 : Umsx84);
	assign G75x84 = (Zapx84 ? Otbw84 : Umsx84);
	assign A75x84 = (Gbpx84 ? Ggdw84 : Umsx84);
	assign U65x84 = (Eapx84 ? Sllw84 : Umsx84);
	assign O65x84 = (X9px84 ? K8nw84 : Umsx84);
	assign I65x84 = (Q9px84 ? Cvow84 : Umsx84);
	assign C65x84 = (J9px84 ? Uhqw84 : Umsx84);
	assign W55x84 = (Nbpx84 ? Y2fw84 : Umsx84);
	assign Q55x84 = (Ubpx84 ? Qpgw84 : Umsx84);
	assign K55x84 = (Bcpx84 ? Iciw84 : Umsx84);
	assign E55x84 = (Icpx84 ? Azjw84 : Umsx84);
	assign Y45x84 = (C9px84 ? M4sw84 : Umsx84);
	assign S45x84 = (V8px84 ? Wdvw84 : Umsx84);
	assign M45x84 = (X4gx84 ? O0xw84 : Umsx84);
	assign Umsx84 = (~(Bnsx84 & Insx84));
	assign Insx84 = (Pnsx84 & Wnsx84);
	assign Wnsx84 = (~(Dosx84 & Uxax84));
	assign Dosx84 = (Ag63a4 & Jgpx84);
	assign Pnsx84 = (Kosx84 & Kdpx84);
	assign Bnsx84 = (Rosx84 & Azjx84);
	assign Azjx84 = (Yosx84 & Fpsx84);
	assign Fpsx84 = (Mpsx84 & Tpsx84);
	assign Tpsx84 = (Aqsx84 | Luqx84);
	assign Mpsx84 = (Hqsx84 & Oqsx84);
	assign Oqsx84 = (Vyrx84 | Ctqx84);
	assign Hqsx84 = (Vqsx84 | Suqx84);
	assign Yosx84 = (Crsx84 & Jrsx84);
	assign Jrsx84 = (Qrsx84 | Qtqx84);
	assign Rosx84 = (Xrsx84 & Essx84);
	assign Essx84 = (~(Qp63a4[25] & Rdpx84));
	assign Xrsx84 = (Shpx84 | Lssx84);
	assign G45x84 = (Gjhx84 ? Attw84 : Sssx84);
	assign A45x84 = (Lapx84 ? Enyw84 : Sssx84);
	assign U35x84 = (Sapx84 ? G60x84 : Sssx84);
	assign O35x84 = (Zapx84 ? Kvbw84 : Sssx84);
	assign I35x84 = (Gbpx84 ? Cidw84 : Sssx84);
	assign C35x84 = (Eapx84 ? Onlw84 : Sssx84);
	assign W25x84 = (X9px84 ? Ganw84 : Sssx84);
	assign Q25x84 = (Q9px84 ? Ywow84 : Sssx84);
	assign K25x84 = (J9px84 ? Qjqw84 : Sssx84);
	assign E25x84 = (Nbpx84 ? U4fw84 : Sssx84);
	assign Y15x84 = (Ubpx84 ? Mrgw84 : Sssx84);
	assign S15x84 = (Bcpx84 ? Eeiw84 : Sssx84);
	assign M15x84 = (Icpx84 ? W0kw84 : Sssx84);
	assign G15x84 = (C9px84 ? I6sw84 : Sssx84);
	assign A15x84 = (V8px84 ? Sfvw84 : Sssx84);
	assign U05x84 = (X4gx84 ? K2xw84 : Sssx84);
	assign Sssx84 = (~(Zssx84 & Gtsx84));
	assign Gtsx84 = (Ntsx84 & Utsx84);
	assign Utsx84 = (~(Busx84 & Nxax84));
	assign Busx84 = (~(Iusx84 | Pusx84));
	assign Ntsx84 = (Wusx84 & Kdpx84);
	assign Zssx84 = (Dvsx84 & Sfkx84);
	assign Sfkx84 = (Kvsx84 & Rvsx84);
	assign Rvsx84 = (Yvsx84 & Fwsx84);
	assign Fwsx84 = (Aqsx84 | J0rx84);
	assign Yvsx84 = (Mwsx84 & Twsx84);
	assign Twsx84 = (Vyrx84 | Ozqx84);
	assign Mwsx84 = (Q0rx84 | Vqsx84);
	assign Kvsx84 = (Crsx84 & Axsx84);
	assign Axsx84 = (Hzqx84 | Qrsx84);
	assign Dvsx84 = (Hxsx84 & Oxsx84);
	assign Oxsx84 = (~(Qp63a4[26] & Rdpx84));
	assign Hxsx84 = (Shpx84 | Vxsx84);
	assign O05x84 = (Gjhx84 ? Wutw84 : Cysx84);
	assign I05x84 = (Lapx84 ? Apyw84 : Cysx84);
	assign Lapx84 = (!Jysx84);
	assign C05x84 = (Sapx84 ? C80x84 : Cysx84);
	assign Sapx84 = (!Qysx84);
	assign Wz4x84 = (Zapx84 ? Gxbw84 : Cysx84);
	assign Zapx84 = (!Xysx84);
	assign Qz4x84 = (Gbpx84 ? Yjdw84 : Cysx84);
	assign Kz4x84 = (Eapx84 ? Kplw84 : Cysx84);
	assign Eapx84 = (!Ezsx84);
	assign Ez4x84 = (X9px84 ? Ccnw84 : Cysx84);
	assign X9px84 = (!Lzsx84);
	assign Yy4x84 = (Q9px84 ? Uyow84 : Cysx84);
	assign Q9px84 = (!Szsx84);
	assign Sy4x84 = (J9px84 ? Mlqw84 : Cysx84);
	assign J9px84 = (!Zzsx84);
	assign My4x84 = (Nbpx84 ? Q6fw84 : Cysx84);
	assign Nbpx84 = (!G0tx84);
	assign Gy4x84 = (Ubpx84 ? Itgw84 : Cysx84);
	assign Ubpx84 = (!N0tx84);
	assign Ay4x84 = (Bcpx84 ? Agiw84 : Cysx84);
	assign Bcpx84 = (!U0tx84);
	assign Ux4x84 = (Icpx84 ? S2kw84 : Cysx84);
	assign Icpx84 = (!B1tx84);
	assign Ox4x84 = (C9px84 ? E8sw84 : Cysx84);
	assign C9px84 = (!I1tx84);
	assign Ix4x84 = (V8px84 ? Ohvw84 : Cysx84);
	assign V8px84 = (!P1tx84);
	assign Cx4x84 = (X4gx84 ? G4xw84 : Cysx84);
	assign Cysx84 = (~(W1tx84 & D2tx84));
	assign D2tx84 = (K2tx84 & R2tx84);
	assign R2tx84 = (~(Y2tx84 & Gxax84));
	assign Y2tx84 = (Hg63a4 & Jgpx84);
	assign K2tx84 = (F3tx84 & Kdpx84);
	assign W1tx84 = (M3tx84 & Cupx84);
	assign Cupx84 = (T3tx84 & A4tx84);
	assign A4tx84 = (H4tx84 & O4tx84);
	assign O4tx84 = (Aqsx84 | M5rx84);
	assign H4tx84 = (V4tx84 & C5tx84);
	assign C5tx84 = (Vyrx84 | R4rx84);
	assign V4tx84 = (T5rx84 | Vqsx84);
	assign T3tx84 = (Crsx84 & J5tx84);
	assign J5tx84 = (K4rx84 | Qrsx84);
	assign M3tx84 = (Q5tx84 & X5tx84);
	assign X5tx84 = (~(Qp63a4[27] & Rdpx84));
	assign Q5tx84 = (Shpx84 | E6tx84);
	assign Ww4x84 = (Gjhx84 ? Swtw84 : L6tx84);
	assign Qw4x84 = (~(S6tx84 & Z6tx84));
	assign Z6tx84 = (G7tx84 | N7tx84);
	assign S6tx84 = (HREADY ? B8tx84 : U7tx84);
	assign B8tx84 = (I8tx84 & P8tx84);
	assign P8tx84 = (~(Wvdx84 & W8tx84));
	assign I8tx84 = (D9tx84 & K9tx84);
	assign K9tx84 = (~(R9tx84 & Y9tx84));
	assign Y9tx84 = (Fatx84 & Matx84);
	assign Fatx84 = (Gv8w84 | Qp63a4[31]);
	assign R9tx84 = (~(Tatx84 | N7tx84));
	assign Tatx84 = (Gqax84 ? Qp63a4[31] : Gv8w84);
	assign D9tx84 = (Mxdx84 | Sgqx84);
	assign U7tx84 = (!Om5w84);
	assign Kw4x84 = (~(Abtx84 & Hbtx84));
	assign Hbtx84 = (Obtx84 & Vbtx84);
	assign Vbtx84 = (~(Czdx84 & Om5w84));
	assign Obtx84 = (~(Jzdx84 & HADDR[28]));
	assign Abtx84 = (Cctx84 & Jctx84);
	assign Jctx84 = (~(E0ex84 & Tk63a4[27]));
	assign Cctx84 = (~(Kcaw84 & L0ex84));
	assign Ew4x84 = (Jysx84 ? L6tx84 : Wqyw84);
	assign Yv4x84 = (Qysx84 ? L6tx84 : Y90x84);
	assign Sv4x84 = (Xysx84 ? L6tx84 : Czbw84);
	assign Mv4x84 = (Gbpx84 ? Uldw84 : L6tx84);
	assign Gv4x84 = (Ezsx84 ? L6tx84 : Grlw84);
	assign Av4x84 = (Lzsx84 ? L6tx84 : Ydnw84);
	assign Uu4x84 = (Szsx84 ? L6tx84 : Q0pw84);
	assign Ou4x84 = (Zzsx84 ? L6tx84 : Inqw84);
	assign Iu4x84 = (G0tx84 ? L6tx84 : M8fw84);
	assign Cu4x84 = (N0tx84 ? L6tx84 : Evgw84);
	assign Wt4x84 = (U0tx84 ? L6tx84 : Whiw84);
	assign Qt4x84 = (B1tx84 ? L6tx84 : O4kw84);
	assign Kt4x84 = (I1tx84 ? L6tx84 : Aasw84);
	assign Et4x84 = (P1tx84 ? L6tx84 : Kjvw84);
	assign Ys4x84 = (X4gx84 ? C6xw84 : L6tx84);
	assign L6tx84 = (~(Qctx84 & Xctx84));
	assign Xctx84 = (Edtx84 & Ldtx84);
	assign Ldtx84 = (~(Qp63a4[28] & Rdpx84));
	assign Edtx84 = (~(Sdtx84 & W8tx84));
	assign Qctx84 = (Sgqx84 & Zdtx84);
	assign Sgqx84 = (Getx84 & Netx84);
	assign Netx84 = (Uetx84 & Bftx84);
	assign Bftx84 = (Aqsx84 | G9rx84);
	assign Uetx84 = (Iftx84 & Pftx84);
	assign Pftx84 = (Vyrx84 | L8rx84);
	assign Iftx84 = (N9rx84 | Vqsx84);
	assign Getx84 = (Crsx84 & Wftx84);
	assign Wftx84 = (E8rx84 | Qrsx84);
	assign Ss4x84 = (Gjhx84 ? Oytw84 : Dgtx84);
	assign Gjhx84 = (!Kgtx84);
	assign Ms4x84 = (~(Rgtx84 & Ygtx84));
	assign Ygtx84 = (~(Th5w84 & Fhtx84));
	assign Fhtx84 = (~(HREADY & Mhtx84));
	assign Mhtx84 = (N7tx84 | Thtx84);
	assign Rgtx84 = (~(HREADY & Aitx84));
	assign Aitx84 = (~(Hitx84 & Oitx84));
	assign Oitx84 = (~(Wvdx84 & Vitx84));
	assign Hitx84 = (Cjtx84 & Jjtx84);
	assign Jjtx84 = (~(Qjtx84 & Ywdx84));
	assign Qjtx84 = (Xjtx84 & Thtx84);
	assign Cjtx84 = (Mxdx84 | Lihx84);
	assign Mxdx84 = (!Ektx84);
	assign Gs4x84 = (~(Lktx84 & Sktx84));
	assign Sktx84 = (Zktx84 & Gltx84);
	assign Gltx84 = (~(Czdx84 & Th5w84));
	assign Zktx84 = (~(Jzdx84 & HADDR[29]));
	assign Lktx84 = (Nltx84 & Ultx84);
	assign Ultx84 = (~(E0ex84 & Tk63a4[28]));
	assign Nltx84 = (~(Geaw84 & L0ex84));
	assign As4x84 = (Jysx84 ? Dgtx84 : Ssyw84);
	assign Ur4x84 = (Qysx84 ? Dgtx84 : Ub0x84);
	assign Or4x84 = (Xysx84 ? Dgtx84 : Y0cw84);
	assign Ir4x84 = (Gbpx84 ? Qndw84 : Dgtx84);
	assign Cr4x84 = (Ezsx84 ? Dgtx84 : Ctlw84);
	assign Wq4x84 = (Lzsx84 ? Dgtx84 : Ufnw84);
	assign Qq4x84 = (Szsx84 ? Dgtx84 : M2pw84);
	assign Kq4x84 = (Zzsx84 ? Dgtx84 : Epqw84);
	assign Eq4x84 = (G0tx84 ? Dgtx84 : Iafw84);
	assign Yp4x84 = (N0tx84 ? Dgtx84 : Axgw84);
	assign Sp4x84 = (U0tx84 ? Dgtx84 : Sjiw84);
	assign Mp4x84 = (B1tx84 ? Dgtx84 : K6kw84);
	assign Gp4x84 = (I1tx84 ? Dgtx84 : Wbsw84);
	assign Ap4x84 = (P1tx84 ? Dgtx84 : Glvw84);
	assign Uo4x84 = (X4gx84 ? Y7xw84 : Dgtx84);
	assign Dgtx84 = (~(Lihx84 & Bmtx84));
	assign Lihx84 = (Imtx84 & Pmtx84);
	assign Pmtx84 = (Wmtx84 & Dntx84);
	assign Dntx84 = (Aqsx84 | Qerx84);
	assign Wmtx84 = (Kntx84 & Rntx84);
	assign Rntx84 = (Vyrx84 | Vdrx84);
	assign Kntx84 = (Xerx84 | Vqsx84);
	assign Imtx84 = (Crsx84 & Yntx84);
	assign Yntx84 = (Odrx84 | Qrsx84);
	assign Oo4x84 = (Kgtx84 ? Q4gx84 : K0uw84);
	assign Q4gx84 = (~(Txdx84 & Fotx84));
	assign Txdx84 = (Motx84 & Totx84);
	assign Totx84 = (Aptx84 & Hptx84);
	assign Hptx84 = (Vyrx84 | Yypx84);
	assign Yypx84 = (Optx84 & Vptx84);
	assign Vptx84 = (Cqtx84 & Jqtx84);
	assign Jqtx84 = (Qqtx84 & Xqtx84);
	assign Xqtx84 = (Ertx84 | Lrtx84);
	assign Qqtx84 = (Srtx84 & Zrtx84);
	assign Srtx84 = (~(Djjx84 & Gstx84));
	assign Cqtx84 = (Nstx84 & Ustx84);
	assign Ustx84 = (~(Bttx84 & Ittx84));
	assign Nstx84 = (~(Pu63a4[14] & Pttx84));
	assign Optx84 = (Wttx84 & Dutx84);
	assign Dutx84 = (Kutx84 & Rutx84);
	assign Rutx84 = (~(X473a4[14] & Yutx84));
	assign Kutx84 = (~(HRDATA[14] & Fvtx84));
	assign Wttx84 = (Mvtx84 & Tvtx84);
	assign Tvtx84 = (~(Nz63a4[2] & Awtx84));
	assign Mvtx84 = (~(STCALIB[14] & Hwtx84));
	assign Aptx84 = (Owtx84 & Vwtx84);
	assign Vwtx84 = (A0qx84 | Vqsx84);
	assign A0qx84 = (Cxtx84 & Jxtx84);
	assign Jxtx84 = (Qxtx84 & Xxtx84);
	assign Xxtx84 = (Eytx84 & Lytx84);
	assign Lytx84 = (~(Bttx84 & Sytx84));
	assign Eytx84 = (Ertx84 | Zytx84);
	assign Qxtx84 = (Gztx84 & Nztx84);
	assign Nztx84 = (~(Pu63a4[22] & Pttx84));
	assign Gztx84 = (~(X473a4[22] & Yutx84));
	assign Cxtx84 = (Uztx84 & B0ux84);
	assign B0ux84 = (I0ux84 & P0ux84);
	assign P0ux84 = (~(HRDATA[22] & Fvtx84));
	assign I0ux84 = (~(W0ux84 & Hw63a4[0]));
	assign Uztx84 = (D1ux84 & K1ux84);
	assign K1ux84 = (~(Nz63a4[4] & Awtx84));
	assign D1ux84 = (~(STCALIB[22] & Hwtx84));
	assign Owtx84 = (Aqsx84 | O0qx84);
	assign O0qx84 = (R1ux84 & Y1ux84);
	assign Y1ux84 = (F2ux84 & M2ux84);
	assign F2ux84 = (T2ux84 & A3ux84);
	assign A3ux84 = (~(H3ux84 & Cahx84));
	assign H3ux84 = (Xx63a4[0] & O3ux84);
	assign T2ux84 = (~(V3ux84 & C4ux84));
	assign R1ux84 = (J4ux84 & Q4ux84);
	assign Q4ux84 = (X4ux84 & E5ux84);
	assign E5ux84 = (~(HRDATA[30] & Fvtx84));
	assign X4ux84 = (~(W0ux84 & D373a4[0]));
	assign J4ux84 = (L5ux84 & S5ux84);
	assign S5ux84 = (~(Nz63a4[6] & Awtx84));
	assign L5ux84 = (~(STCALIB[24] & Hwtx84));
	assign Motx84 = (Crsx84 & Z5ux84);
	assign Z5ux84 = (Q1qx84 | Qrsx84);
	assign Q1qx84 = (G6ux84 & N6ux84);
	assign N6ux84 = (U6ux84 & B7ux84);
	assign B7ux84 = (I7ux84 & P7ux84);
	assign P7ux84 = (~(Bttx84 & W7ux84));
	assign I7ux84 = (Ertx84 | D8ux84);
	assign U6ux84 = (K8ux84 & R8ux84);
	assign R8ux84 = (~(Pu63a4[6] & Pttx84));
	assign K8ux84 = (~(X473a4[6] & Yutx84));
	assign G6ux84 = (Y8ux84 & F9ux84);
	assign F9ux84 = (~(STCALIB[6] & Hwtx84));
	assign Y8ux84 = (M9ux84 & T9ux84);
	assign T9ux84 = (~(HRDATA[6] & Fvtx84));
	assign M9ux84 = (~(Nz63a4[0] & Awtx84));
	assign Io4x84 = (Kgtx84 ? E5gx84 : G2uw84);
	assign E5gx84 = (Mqdx84 | Aaux84);
	assign Co4x84 = (~(Haux84 & Oaux84));
	assign Oaux84 = (Vaux84 & Cbux84);
	assign Cbux84 = (~(Cr63a4[15] & Hrdx84));
	assign Vaux84 = (Jbux84 & Qbux84);
	assign Qbux84 = (Igex84 | Xbux84);
	assign Jbux84 = (~(Qp63a4[16] & Kpdx84));
	assign Haux84 = (Jbgx84 & Ecux84);
	assign Ecux84 = (~(Tk63a4[15] & Ordx84));
	assign Jbgx84 = (Lcux84 & Ypdx84);
	assign Lcux84 = (Igex84 | Czrx84);
	assign Wn4x84 = (Jysx84 ? Scux84 : S4yw84);
	assign Qn4x84 = (Qysx84 ? Scux84 : Unzw84);
	assign Kn4x84 = (Xysx84 ? Scux84 : Ycbw84);
	assign En4x84 = (Gbpx84 ? Qzcw84 : Scux84);
	assign Ym4x84 = (Ezsx84 ? Scux84 : C5lw84);
	assign Sm4x84 = (Lzsx84 ? Scux84 : Urmw84);
	assign Mm4x84 = (Szsx84 ? Scux84 : Meow84);
	assign Gm4x84 = (Zzsx84 ? Scux84 : E1qw84);
	assign Am4x84 = (G0tx84 ? Scux84 : Imew84);
	assign Ul4x84 = (N0tx84 ? Scux84 : A9gw84);
	assign Ol4x84 = (U0tx84 ? Scux84 : Svhw84);
	assign Il4x84 = (B1tx84 ? Scux84 : Kijw84);
	assign Cl4x84 = (I1tx84 ? Scux84 : Wnrw84);
	assign Wk4x84 = (Kgtx84 ? Scux84 : Oatw84);
	assign Qk4x84 = (P1tx84 ? Scux84 : Gxuw84);
	assign Kk4x84 = (X4gx84 ? Yjww84 : Scux84);
	assign Scux84 = (~(Zcux84 & Gdux84));
	assign Gdux84 = (Ndux84 & Udux84);
	assign Udux84 = (~(Qp63a4[16] & Rdpx84));
	assign Ndux84 = (Beux84 & Ieux84);
	assign Beux84 = (~(Peux84 & M0bx84));
	assign Peux84 = (Jgpx84 & Ch63a4);
	assign Jgpx84 = (!Iusx84);
	assign Zcux84 = (Weux84 & Xbux84);
	assign Xbux84 = (Dfux84 & Kfux84);
	assign Kfux84 = (Rfux84 & Yfux84);
	assign Yfux84 = (Mxrx84 | Bpqx84);
	assign Mxrx84 = (Qsrx84 & Unrx84);
	assign Rfux84 = (Txrx84 | Dqqx84);
	assign Txrx84 = (Rprx84 ? Fgux84 : Raex84);
	assign Dfux84 = (Mgux84 & Tgux84);
	assign Tgux84 = (Oyrx84 | Rqqx84);
	assign Oyrx84 = (Ahux84 | Hhux84);
	assign Mgux84 = (Vyrx84 | Noqx84);
	assign Weux84 = (N8sx84 & Ohux84);
	assign Ohux84 = (Shpx84 | Vhux84);
	assign N8sx84 = (Czrx84 & Kdpx84);
	assign Czrx84 = (Ciux84 & Jiux84);
	assign Ciux84 = (~(Qiux84 & Hhux84));
	assign Qiux84 = (Xiux84 & Fgux84);
	assign Ek4x84 = (~(Ejux84 & Ljux84));
	assign Ljux84 = (Sjux84 & Zjux84);
	assign Zjux84 = (~(Kpdx84 & Qp63a4[24]));
	assign Kpdx84 = (Izgx84 & R3ex84);
	assign Sjux84 = (Gkux84 & Ypdx84);
	assign Ypdx84 = (~(Izgx84 & Nkux84));
	assign Nkux84 = (~(Ukux84 & Blux84));
	assign Blux84 = (~(Nx4w84 & Ilux84));
	assign Ukux84 = (Plux84 & W2ex84);
	assign W2ex84 = (!LOCKUP);
	assign Plux84 = (~(Wlux84 & Uv4w84));
	assign Wlux84 = (Nj63a4[0] & Dmux84);
	assign Gkux84 = (Igex84 | M4ex84);
	assign Igex84 = (!Fqdx84);
	assign Fqdx84 = (~(T4ex84 | Ordx84));
	assign Ejux84 = (Kmux84 & Rmux84);
	assign Rmux84 = (~(Cr63a4[23] & Hrdx84));
	assign Hrdx84 = (Ymux84 & Fnux84);
	assign Ymux84 = (Izgx84 & T4ex84);
	assign T4ex84 = (!Soix84);
	assign Kmux84 = (~(Tk63a4[23] & Ordx84));
	assign Ordx84 = (!Izgx84);
	assign Izgx84 = (HREADY & Mnux84);
	assign Yj4x84 = (~(Tnux84 & Aoux84));
	assign Aoux84 = (Houx84 & Ooux84);
	assign Ooux84 = (~(P25w84 & Czdx84));
	assign Houx84 = (~(Jzdx84 & HADDR[24]));
	assign Tnux84 = (Voux84 & Cpux84);
	assign Cpux84 = (~(Tk63a4[23] & E0ex84));
	assign Voux84 = (~(A5aw84 & L0ex84));
	assign Sj4x84 = (Jysx84 ? Jpux84 : Mjyw84);
	assign Jysx84 = (Qpux84 & Xpux84);
	assign Qpux84 = (~(Fvfx84 | Equx84));
	assign Mj4x84 = (Qysx84 ? Jpux84 : O20x84);
	assign Qysx84 = (Lqux84 & Xpux84);
	assign Lqux84 = (~(Equx84 | Mdxw84));
	assign Gj4x84 = (Xysx84 ? Jpux84 : Srbw84);
	assign Xysx84 = (Squx84 & Zqux84);
	assign Squx84 = (~(Grux84 | Nrux84));
	assign Aj4x84 = (Gbpx84 ? Kedw84 : Jpux84);
	assign Gbpx84 = (~(Xpux84 & Equx84));
	assign Xpux84 = (Urux84 & Bsux84);
	assign Urux84 = (Isux84 & Psux84);
	assign Ui4x84 = (Ezsx84 ? Jpux84 : Wjlw84);
	assign Ezsx84 = (Wsux84 & Dtux84);
	assign Wsux84 = (~(Psux84 | Nrux84));
	assign Oi4x84 = (Lzsx84 ? Jpux84 : O6nw84);
	assign Lzsx84 = (Ktux84 & Rtux84);
	assign Ktux84 = (~(Nrux84 | Bsux84));
	assign Ii4x84 = (Szsx84 ? Jpux84 : Gtow84);
	assign Szsx84 = (Ytux84 & Fuux84);
	assign Fuux84 = (~(Nrux84 | Equx84));
	assign Ytux84 = (~(Muux84 | Psux84));
	assign Ci4x84 = (Zzsx84 ? Jpux84 : Yfqw84);
	assign Zzsx84 = (Tuux84 & Rtux84);
	assign Tuux84 = (~(Muux84 | Nrux84));
	assign Nrux84 = (!Isux84);
	assign Wh4x84 = (G0tx84 ? Jpux84 : C1fw84);
	assign G0tx84 = (Avux84 & Hvux84);
	assign Qh4x84 = (N0tx84 ? Jpux84 : Ungw84);
	assign N0tx84 = (Ovux84 & Zqux84);
	assign Zqux84 = (Muux84 & Psux84);
	assign Ovux84 = (~(Isux84 | Grux84));
	assign Kh4x84 = (U0tx84 ? Jpux84 : Maiw84);
	assign U0tx84 = (Hvux84 & Vvux84);
	assign Hvux84 = (Grux84 & Psux84);
	assign Eh4x84 = (B1tx84 ? Jpux84 : Exjw84);
	assign B1tx84 = (Cwux84 & Vvux84);
	assign Cwux84 = (Equx84 & Psux84);
	assign Yg4x84 = (I1tx84 ? Jpux84 : Q2sw84);
	assign I1tx84 = (Jwux84 & Dtux84);
	assign Dtux84 = (~(Bsux84 | Equx84));
	assign Jwux84 = (~(Isux84 | Psux84));
	assign Sg4x84 = (Kgtx84 ? Jpux84 : Iptw84);
	assign Kgtx84 = (Avux84 & Rtux84);
	assign Avux84 = (~(Isux84 | Bsux84));
	assign Bsux84 = (!Muux84);
	assign Mg4x84 = (P1tx84 ? Jpux84 : Acvw84);
	assign P1tx84 = (Qwux84 & Vvux84);
	assign Qwux84 = (~(Psux84 | Equx84));
	assign Equx84 = (!Grux84);
	assign Gg4x84 = (X4gx84 ? Syww84 : Jpux84);
	assign X4gx84 = (~(Rtux84 & Vvux84));
	assign Vvux84 = (~(Muux84 | Isux84));
	assign Isux84 = (~(Xwux84 & Exux84));
	assign Exux84 = (Lxux84 & Sxux84);
	assign Sxux84 = (Zxux84 | Gyux84);
	assign Lxux84 = (Nyux84 & Uyux84);
	assign Uyux84 = (Bzux84 | Izux84);
	assign Nyux84 = (Tmox84 | Pzux84);
	assign Muux84 = (~(Wzux84 & D0vx84));
	assign D0vx84 = (K0vx84 & HREADY);
	assign K0vx84 = (R0vx84 & Y0vx84);
	assign Wzux84 = (F1vx84 & M1vx84);
	assign Rtux84 = (~(Psux84 | Grux84));
	assign Grux84 = (~(T1vx84 & A2vx84));
	assign A2vx84 = (H2vx84 & O2vx84);
	assign O2vx84 = (V2vx84 | Izux84);
	assign H2vx84 = (Dnmx84 | Pzux84);
	assign T1vx84 = (C3vx84 & J3vx84);
	assign J3vx84 = (Q3vx84 | Gyux84);
	assign Psux84 = (~(Xwux84 & X3vx84));
	assign X3vx84 = (E4vx84 & L4vx84);
	assign L4vx84 = (S4vx84 | Gyux84);
	assign E4vx84 = (Z4vx84 & G5vx84);
	assign G5vx84 = (N5vx84 | Izux84);
	assign Z4vx84 = (T7px84 | Pzux84);
	assign Xwux84 = (C3vx84 & M1vx84);
	assign C3vx84 = (U5vx84 & HREADY);
	assign U5vx84 = (B6vx84 & R0vx84);
	assign R0vx84 = (~(I6vx84 & P6vx84));
	assign P6vx84 = (W6vx84 & D7vx84);
	assign D7vx84 = (K7vx84 & R7vx84);
	assign R7vx84 = (~(Hghx84 & Y7vx84));
	assign Y7vx84 = (~(F8vx84 & M8vx84));
	assign M8vx84 = (~(T8vx84 & N4ix84));
	assign T8vx84 = (~(Evix84 | Zo2x84));
	assign F8vx84 = (O8bx84 | Gpbx84);
	assign K7vx84 = (A9vx84 & H9vx84);
	assign H9vx84 = (~(O9vx84 & Phdx84));
	assign O9vx84 = (~(F5dx84 | Yqcx84));
	assign A9vx84 = (~(Atix84 & V9vx84));
	assign V9vx84 = (Cavx84 | Javx84);
	assign W6vx84 = (Qavx84 & Xavx84);
	assign Xavx84 = (~(Krix84 & T0px84));
	assign Qavx84 = (Ebvx84 & Lbvx84);
	assign Lbvx84 = (~(Sbvx84 & Zbvx84));
	assign Zbvx84 = (Jsrx84 | T0px84);
	assign Ebvx84 = (~(Gcvx84 & Ncvx84));
	assign Ncvx84 = (~(Wtfx84 & Ucvx84));
	assign Ucvx84 = (Gzfx84 | J13x84);
	assign I6vx84 = (Bdvx84 & Idvx84);
	assign Idvx84 = (Pdvx84 & Wdvx84);
	assign Wdvx84 = (~(E3ix84 & Devx84));
	assign Pdvx84 = (Kevx84 & Revx84);
	assign Revx84 = (~(Yevx84 & Hbmx84));
	assign Kevx84 = (~(Vx2x84 & Ffvx84));
	assign Ffvx84 = (~(Mfvx84 & Tfvx84));
	assign Tfvx84 = (~(Agvx84 & Hgvx84));
	assign Agvx84 = (Ogvx84 | Vgvx84);
	assign Vgvx84 = (Dzox84 & H6dx84);
	assign Mfvx84 = (Chvx84 & Jhvx84);
	assign Jhvx84 = (~(Qhvx84 & Xhvx84));
	assign Qhvx84 = (~(Jnix84 | J13x84));
	assign Chvx84 = (~(Eivx84 & Livx84));
	assign Eivx84 = (~(Yqcx84 | Pqbx84));
	assign Bdvx84 = (Sivx84 & Zivx84);
	assign Zivx84 = (Pqbx84 ? Njvx84 : Gjvx84);
	assign Njvx84 = (Ujvx84 & Bkvx84);
	assign Bkvx84 = (Ikvx84 & P1mx84);
	assign Ikvx84 = (~(Pkvx84 & Gz4w84));
	assign Pkvx84 = (~(Hu2x84 | Bw2x84));
	assign Ujvx84 = (Wkvx84 & Dlvx84);
	assign Dlvx84 = (~(Yevx84 & Klvx84));
	assign Wkvx84 = (Fn2x84 | J13x84);
	assign Sivx84 = (Rlvx84 & Ylvx84);
	assign Rlvx84 = (B0gx84 | H6dx84);
	assign B6vx84 = (Fmvx84 | Mmvx84);
	assign Jpux84 = (~(M4ex84 & Tmvx84));
	assign M4ex84 = (Anvx84 & Hnvx84);
	assign Hnvx84 = (Onvx84 & Vnvx84);
	assign Vnvx84 = (Aqsx84 | Dqqx84);
	assign Onvx84 = (Covx84 & Jovx84);
	assign Jovx84 = (Vyrx84 | Bpqx84);
	assign Covx84 = (Rqqx84 | Vqsx84);
	assign Anvx84 = (Crsx84 & Qovx84);
	assign Qovx84 = (Noqx84 | Qrsx84);
	assign Ag4x84 = (~(Xovx84 & Epvx84));
	assign Epvx84 = (Lpvx84 & Spvx84);
	assign Spvx84 = (~(Zpvx84 & Gqvx84));
	assign Gqvx84 = (~(Nqvx84 | Shix84));
	assign Zpvx84 = (Jzdx84 & Uqvx84);
	assign Uqvx84 = (Gpbx84 | Gf6w84);
	assign Lpvx84 = (~(Czdx84 & Nj63a4[1]));
	assign Xovx84 = (Brvx84 & Irvx84);
	assign Irvx84 = (~(E0ex84 & Tk63a4[0]));
	assign Brvx84 = (~(Xy8w84 & L0ex84));
	assign Uf4x84 = (Bvdx84 ? Prvx84 : Up5w84);
	assign Bvdx84 = (HREADY & Wrvx84);
	assign Wrvx84 = (N7tx84 | Dsvx84);
	assign N7tx84 = (!Ywdx84);
	assign Prvx84 = (~(Ksvx84 & Rsvx84));
	assign Rsvx84 = (~(Wvdx84 & Ysvx84));
	assign Ksvx84 = (Ftvx84 & Mtvx84);
	assign Mtvx84 = (~(Ttvx84 & Ywdx84));
	assign Ywdx84 = (~(Wvdx84 | Ektx84));
	assign Wvdx84 = (Auvx84 & P7gx84);
	assign Ftvx84 = (~(Ektx84 & Mqdx84));
	assign Mqdx84 = (~(Huvx84 & Ouvx84));
	assign Ouvx84 = (Vuvx84 & Cvvx84);
	assign Cvvx84 = (Aqsx84 | Hlqx84);
	assign Aqsx84 = (Jvvx84 | Ahux84);
	assign Ahux84 = (Qvvx84 & Gz4w84);
	assign Qvvx84 = (~(Rprx84 | Deox84));
	assign Vuvx84 = (Xvvx84 & Ewvx84);
	assign Ewvx84 = (Vyrx84 | Olqx84);
	assign Vyrx84 = (~(Lwvx84 & Rprx84));
	assign Xvvx84 = (Vqsx84 | Cmqx84);
	assign Vqsx84 = (Unrx84 & Swvx84);
	assign Swvx84 = (Raex84 | Rprx84);
	assign Unrx84 = (Zwvx84 | Orrx84);
	assign Huvx84 = (Crsx84 & Gxvx84);
	assign Gxvx84 = (Qrsx84 | Mkqx84);
	assign Qrsx84 = (Qsrx84 & Nxvx84);
	assign Nxvx84 = (Uxvx84 | Orrx84);
	assign Crsx84 = (Byvx84 & Jiux84);
	assign Jiux84 = (~(Iyvx84 & Pyvx84));
	assign Pyvx84 = (~(Wyvx84 & Dzvx84));
	assign Dzvx84 = (~(P0gx84 & Mmvx84));
	assign Wyvx84 = (Kzvx84 & Pvrx84);
	assign Iyvx84 = (Gurx84 & Orrx84);
	assign Byvx84 = (~(Rzvx84 & Xiux84));
	assign Xiux84 = (Yzvx84 & F0wx84);
	assign Yzvx84 = (Gurx84 & Zwvx84);
	assign Rzvx84 = (Jvvx84 & Uxvx84);
	assign Jvvx84 = (Rprx84 & M0wx84);
	assign Ektx84 = (T0wx84 & Hscx84);
	assign Of4x84 = (Eabx84 ? A1wx84 : Iv6w84);
	assign Eabx84 = (HREADY & H1wx84);
	assign H1wx84 = (~(O1wx84 & V1wx84));
	assign V1wx84 = (C2wx84 & J2wx84);
	assign J2wx84 = (Q2wx84 & X2wx84);
	assign X2wx84 = (~(E3wx84 & L3wx84));
	assign L3wx84 = (~(S3wx84 & Z3wx84));
	assign Z3wx84 = (Jxmx84 | G4wx84);
	assign S3wx84 = (N4wx84 & U4wx84);
	assign N4wx84 = (~(B5wx84 & Kprx84));
	assign B5wx84 = (~(Fmvx84 | Vx2x84));
	assign Q2wx84 = (I5wx84 & P5wx84);
	assign I5wx84 = (~(W5wx84 & W05w84));
	assign W5wx84 = (Gpix84 & Gknx84);
	assign Gknx84 = (~(D6wx84 & K6wx84));
	assign K6wx84 = (Fmvx84 | Ewax84);
	assign D6wx84 = (Gz4w84 | Ns2x84);
	assign C2wx84 = (R6wx84 & Y6wx84);
	assign Y6wx84 = (~(Gz4w84 & F7wx84));
	assign F7wx84 = (~(M7wx84 & T7wx84));
	assign T7wx84 = (~(Lzlx84 & A8wx84));
	assign A8wx84 = (~(Efdx84 & H8wx84));
	assign H8wx84 = (~(O8wx84 & V8wx84));
	assign M7wx84 = (~(Uemx84 & Ba6w84));
	assign R6wx84 = (~(S6mx84 & C9wx84));
	assign O1wx84 = (J9wx84 & Q9wx84);
	assign Q9wx84 = (X9wx84 & D2mx84);
	assign D2mx84 = (Eawx84 & Lawx84);
	assign Lawx84 = (Sawx84 & Zawx84);
	assign Zawx84 = (~(Gbwx84 & Nbwx84));
	assign Nbwx84 = (~(Gpbx84 | Lfdx84));
	assign Gbwx84 = (Ubwx84 & C2ix84);
	assign Sawx84 = (~(Benx84 & F3mx84));
	assign Eawx84 = (Aonx84 & Bcwx84);
	assign Bcwx84 = (~(Huhx84 & Zg6w84));
	assign Aonx84 = (Icwx84 & Qxfx84);
	assign Qxfx84 = (Xubx84 | J8cx84);
	assign Icwx84 = (Pcwx84 & Cubx84);
	assign Pcwx84 = (~(Wcwx84 & E9cx84));
	assign X9wx84 = (Ddwx84 & Kdwx84);
	assign Kdwx84 = (Xubx84 | Xlkx84);
	assign Ddwx84 = (Saix84 | Yqcx84);
	assign Saix84 = (!Hbmx84);
	assign J9wx84 = (Bsnx84 & Tnnx84);
	assign Tnnx84 = (Rdwx84 & Ydwx84);
	assign Ydwx84 = (~(L2cx84 & C2ix84));
	assign Rdwx84 = (~(Dzox84 & Gpbx84));
	assign Bsnx84 = (Fewx84 & Mewx84);
	assign Mewx84 = (~(Pxbx84 & Tewx84));
	assign Tewx84 = (~(Afwx84 & Hfwx84));
	assign Hfwx84 = (Fthx84 | Fn2x84);
	assign Afwx84 = (Ofwx84 & Vfwx84);
	assign Ofwx84 = (~(E3wx84 & Laix84));
	assign Fewx84 = (Cgwx84 & Jgwx84);
	assign Jgwx84 = (~(Qgwx84 & Devx84));
	assign Qgwx84 = (Xgwx84 & Wqbx84);
	assign Cgwx84 = (~(Ehwx84 & V1ix84));
	assign Ehwx84 = (~(J8cx84 | Fcdx84));
	assign A1wx84 = (~(Lhwx84 & Shwx84));
	assign Shwx84 = (Zhwx84 & Giwx84);
	assign Giwx84 = (~(Y46w84 & Niwx84));
	assign Niwx84 = (~(Ijbx84 & Rdbx84));
	assign Rdbx84 = (~(Uiwx84 & Fcdx84));
	assign Uiwx84 = (~(I4cx84 | Cfcx84));
	assign Ijbx84 = (Bjwx84 & R7ox84);
	assign R7ox84 = (Ijwx84 & U9dx84);
	assign U9dx84 = (Cfcx84 | Ub6w84);
	assign Ijwx84 = (~(Pjwx84 & Evbx84));
	assign Bjwx84 = (Wjwx84 & Kdbx84);
	assign Kdbx84 = (~(Dkwx84 & Kkwx84));
	assign Kkwx84 = (~(Rkwx84 & Xubx84));
	assign Rkwx84 = (~(Ykwx84 | B9lx84));
	assign Dkwx84 = (E8dx84 | Fhmx84);
	assign Zhwx84 = (~(Kr5w84 & Uibx84));
	assign Uibx84 = (~(Flwx84 & Bcbx84));
	assign Bcbx84 = (Xgix84 & Mlwx84);
	assign Mlwx84 = (~(Tlwx84 & Pcbx84));
	assign Xgix84 = (~(Huhx84 & Edmx84));
	assign Flwx84 = (Amwx84 & Hmwx84);
	assign Hmwx84 = (~(E8dx84 & Omwx84));
	assign Omwx84 = (~(Vmwx84 & Cnwx84));
	assign Cnwx84 = (~(C9wx84 & J8cx84));
	assign C9wx84 = (~(Jnwx84 & E2cx84));
	assign Vmwx84 = (~(Huhx84 & Xlkx84));
	assign Amwx84 = (~(Pcbx84 & Z6mx84));
	assign Lhwx84 = (Ydbx84 & Qnwx84);
	assign Qnwx84 = (Mebx84 | Qzkx84);
	assign Ydbx84 = (Xnwx84 & Eowx84);
	assign Eowx84 = (~(Lowx84 | Zymx84));
	assign Xnwx84 = (Sowx84 & Zowx84);
	assign Zowx84 = (~(Xlkx84 & Gpwx84));
	assign Gpwx84 = (~(Npwx84 & T7ix84));
	assign T7ix84 = (~(Upwx84 & W05w84));
	assign Upwx84 = (~(Bqwx84 | Fn2x84));
	assign Npwx84 = (~(Symx84 | B9lx84));
	assign Sowx84 = (~(Wadx84 & G36w84));
	assign If4x84 = (!Iqwx84);
	assign Iqwx84 = (HREADY ? Pqwx84 : Xvax84);
	assign Pqwx84 = (Wqwx84 & Drwx84);
	assign Drwx84 = (Krwx84 & Rrwx84);
	assign Rrwx84 = (Yrwx84 & Fswx84);
	assign Fswx84 = (~(Mswx84 & Qvax84));
	assign Mswx84 = (~(Tswx84 | Tq2x84));
	assign Yrwx84 = (Atwx84 & Lcnx84);
	assign Lcnx84 = (~(Htwx84 & Nndx84));
	assign Htwx84 = (~(Qxmx84 | Gz4w84));
	assign Atwx84 = (~(Otwx84 & Uwix84));
	assign Otwx84 = (~(Lrfx84 | Wqbx84));
	assign Krwx84 = (Vtwx84 & Cuwx84);
	assign Cuwx84 = (~(Atix84 & Juwx84));
	assign Juwx84 = (Quwx84 | Xuwx84);
	assign Xuwx84 = (W05w84 ? Zg6w84 : Evwx84);
	assign Evwx84 = (~(Lvwx84 & Svwx84));
	assign Svwx84 = (~(Zvwx84 & J8cx84));
	assign Zvwx84 = (Nd6w84 | X8cx84);
	assign Lvwx84 = (~(Uemx84 & Gwwx84));
	assign Gwwx84 = (~(Nwwx84 & Uwwx84));
	assign Uwwx84 = (~(Nrnx84 | Ub6w84));
	assign Nwwx84 = (Bxwx84 & Ixwx84);
	assign Bxwx84 = (Eobx84 ? G36w84 : Pxwx84);
	assign Quwx84 = (~(Wxwx84 & Dywx84));
	assign Dywx84 = (~(Kywx84 & Ybdx84));
	assign Ybdx84 = (Hddx84 ^ Eobx84);
	assign Hddx84 = (~(Rywx84 & Yywx84));
	assign Yywx84 = (Fzwx84 ^ Mzwx84);
	assign Mzwx84 = (~(Tzwx84 | A0xx84));
	assign A0xx84 = (Dsvx84 ? Ttvx84 : Up5w84);
	assign Ttvx84 = (~(H0xx84 | O0xx84));
	assign O0xx84 = (V0xx84 & Me5w84);
	assign Tzwx84 = (Qqmx84 | Ixwx84);
	assign Fzwx84 = (~(C1xx84 & J1xx84));
	assign J1xx84 = (G7tx84 & Q1xx84);
	assign G7tx84 = (~(X1xx84 & Om5w84));
	assign X1xx84 = (E2xx84 & L2xx84);
	assign C1xx84 = (S2xx84 & Bfmx84);
	assign Bfmx84 = (~(Tqkx84 & Z6mx84));
	assign S2xx84 = (~(Z2xx84 & G3xx84));
	assign G3xx84 = (Gqax84 ? Gv8w84 : Qp63a4[31]);
	assign Z2xx84 = (N3xx84 & Matx84);
	assign Matx84 = (~(E2xx84 & L2xx84));
	assign L2xx84 = (~(Pqbx84 & U3xx84));
	assign U3xx84 = (~(B4xx84 & F5dx84));
	assign B4xx84 = (~(Sbvx84 & I4xx84));
	assign I4xx84 = (~(P4xx84 & W4xx84));
	assign W4xx84 = (Wqbx84 | Fn2x84);
	assign P4xx84 = (D5xx84 & K5xx84);
	assign D5xx84 = (Evix84 | Zo2x84);
	assign E2xx84 = (~(Gz4w84 & R5xx84));
	assign R5xx84 = (~(Y5xx84 & F6xx84));
	assign F6xx84 = (M6xx84 | D4dx84);
	assign Y5xx84 = (T6xx84 & A7xx84);
	assign A7xx84 = (~(H7xx84 & Livx84));
	assign H7xx84 = (~(Jnix84 | Zo2x84));
	assign T6xx84 = (Sbox84 | Mmvx84);
	assign N3xx84 = (~(Gv8w84 & Qp63a4[31]));
	assign Gv8w84 = (O7xx84 & Q2bx84);
	assign Q2bx84 = (~(V7xx84 & C8xx84));
	assign C8xx84 = (J8xx84 & Q8xx84);
	assign Q8xx84 = (X8xx84 & E9xx84);
	assign E9xx84 = (~(Pxbx84 & L9xx84));
	assign L9xx84 = (Undx84 | Deox84);
	assign X8xx84 = (~(S9xx84 | Hbmx84));
	assign J8xx84 = (Z9xx84 & Gaxx84);
	assign Gaxx84 = (Naxx84 | B5bx84);
	assign Z9xx84 = (Uaxx84 & Bbxx84);
	assign Bbxx84 = (Zbox84 | Bw2x84);
	assign Uaxx84 = (Xqfx84 | Hu2x84);
	assign V7xx84 = (Ibxx84 & Pbxx84);
	assign Pbxx84 = (Wbxx84 & Dcxx84);
	assign Dcxx84 = (Ewax84 | Evix84);
	assign Wbxx84 = (Ibcx84 & Kcxx84);
	assign Kcxx84 = (Yshx84 | Fycx84);
	assign Ibcx84 = (F5dx84 | G4bx84);
	assign Ibxx84 = (Ol2x84 & Rcxx84);
	assign Rcxx84 = (Pqbx84 | J13x84);
	assign Rywx84 = (Ycxx84 & Fdxx84);
	assign Fdxx84 = (Mdxx84 | Tdxx84);
	assign Tdxx84 = (Thtx84 ? Xjtx84 : Th5w84);
	assign Thtx84 = (~(Aexx84 & Hexx84));
	assign Hexx84 = (Gjvx84 & Oexx84);
	assign Oexx84 = (~(Hghx84 & Nndx84));
	assign Aexx84 = (Vexx84 & Cfxx84);
	assign Cfxx84 = (~(Jfxx84 & F7bx84));
	assign Vexx84 = (~(Pqbx84 & Qfxx84));
	assign Qfxx84 = (~(Xfxx84 & Egxx84));
	assign Egxx84 = (~(Lgxx84 & Yzhx84));
	assign Lgxx84 = (~(Fn2x84 | J13x84));
	assign Xfxx84 = (~(Sbvx84 & Sgxx84));
	assign Sgxx84 = (Zgxx84 | Ghxx84);
	assign Xjtx84 = (Me5w84 ? Nhxx84 : S17w84);
	assign Nhxx84 = (Bixx84 ? Th5w84 : Uhxx84);
	assign Bixx84 = (Iixx84 & Pixx84);
	assign Uhxx84 = (~(Wixx84 & Djxx84));
	assign Djxx84 = (~(Kjxx84 & Rjxx84));
	assign Rjxx84 = (~(Yjxx84 & Wbcx84));
	assign Yjxx84 = (~(Fkxx84 & Mkxx84));
	assign Kjxx84 = (~(Tkxx84 & Alxx84));
	assign Alxx84 = (~(Hlxx84 & Olxx84));
	assign Hlxx84 = (Vlxx84 & Cmxx84);
	assign Tkxx84 = (~(Jmxx84 & Qmxx84));
	assign Qmxx84 = (~(Xmxx84 & Cmxx84));
	assign Jmxx84 = (Olxx84 ? Lnxx84 : Enxx84);
	assign Lnxx84 = (~(Snxx84 | Cmxx84));
	assign Enxx84 = (Cmxx84 | Znxx84);
	assign Wixx84 = (Mkxx84 ? Noxx84 : Goxx84);
	assign Mkxx84 = (Uoxx84 | Iixx84);
	assign Uoxx84 = (Pixx84 & Bpxx84);
	assign Pixx84 = (!Ipxx84);
	assign Noxx84 = (~(Ppxx84 & Wpxx84));
	assign Ppxx84 = (~(Dqxx84 & Kqxx84));
	assign Kqxx84 = (~(Rqxx84 & Yqxx84));
	assign Dqxx84 = (Olxx84 ? Mrxx84 : Frxx84);
	assign Mrxx84 = (!Trxx84);
	assign Trxx84 = (Osxx84 ? Hsxx84 : Asxx84);
	assign Frxx84 = (~(Osxx84 & Vsxx84));
	assign Goxx84 = (Bqwx84 | V0xx84);
	assign V0xx84 = (Ctxx84 & Jtxx84);
	assign Jtxx84 = (Qtxx84 & Xtxx84);
	assign Xtxx84 = (~(Lwvx84 & Vlxx84));
	assign Qtxx84 = (Euxx84 & Luxx84);
	assign Euxx84 = (Uxvx84 | Suxx84);
	assign Ctxx84 = (Zuxx84 & Gvxx84);
	assign Gvxx84 = (Zwvx84 | Snxx84);
	assign Zuxx84 = (~(Nvxx84 & Uvxx84));
	assign Mdxx84 = (~(Bwxx84 & Tebx84));
	assign Bwxx84 = (Qqmx84 | Iwxx84);
	assign Ycxx84 = (~(Pwxx84 & Wwxx84));
	assign Wwxx84 = (Dxxx84 ^ Gwbx84);
	assign Dxxx84 = (Kxxx84 ? Eo5w84 : Fxdx84);
	assign Kxxx84 = (!Dsvx84);
	assign Dsvx84 = (~(Rxxx84 & Yxxx84));
	assign Yxxx84 = (Fyxx84 & Myxx84);
	assign Myxx84 = (~(Tyxx84 & Gz4w84));
	assign Tyxx84 = (~(D4dx84 | Hu2x84));
	assign Fyxx84 = (Azxx84 & Gjvx84);
	assign Gjvx84 = (~(Hzxx84 & Klvx84));
	assign Hzxx84 = (~(F5dx84 | Zo2x84));
	assign Azxx84 = (~(Ozxx84 & F7bx84));
	assign Ozxx84 = (~(F5dx84 | Wqbx84));
	assign Rxxx84 = (Vzxx84 & C0yx84);
	assign C0yx84 = (~(Pqbx84 & J0yx84));
	assign J0yx84 = (Hghx84 | Q0yx84);
	assign Vzxx84 = (~(Nndx84 & Gz4w84));
	assign Fxdx84 = (~(X0yx84 & E1yx84));
	assign E1yx84 = (~(L1yx84 & S1yx84));
	assign S1yx84 = (Z1yx84 & G2yx84);
	assign G2yx84 = (~(N2yx84 & U2yx84));
	assign U2yx84 = (~(B3yx84 & I3yx84));
	assign I3yx84 = (P3yx84 & Zytx84);
	assign P3yx84 = (~(Asxx84 | W3yx84));
	assign W3yx84 = (!Snxx84);
	assign B3yx84 = (D4yx84 & K4yx84);
	assign D4yx84 = (F5yx84 ? Y4yx84 : R4yx84);
	assign Y4yx84 = (M5yx84 & T5yx84);
	assign T5yx84 = (A6yx84 & H6yx84);
	assign M5yx84 = (~(O6yx84 | Sytx84));
	assign R4yx84 = (V6yx84 & C7yx84);
	assign C7yx84 = (~(J7yx84 | Q7yx84));
	assign N2yx84 = (~(X7yx84 & Uurx84));
	assign Z1yx84 = (E8yx84 & Luxx84);
	assign E8yx84 = (~(L8yx84 & S8yx84));
	assign S8yx84 = (~(Z8yx84 & G9yx84));
	assign G9yx84 = (N9yx84 & Lrtx84);
	assign N9yx84 = (~(Vsxx84 | Vlxx84));
	assign Z8yx84 = (U9yx84 & Bayx84);
	assign U9yx84 = (F5yx84 ? Payx84 : Iayx84);
	assign Payx84 = (V6yx84 & Wayx84);
	assign Wayx84 = (~(Dbyx84 | Kbyx84));
	assign V6yx84 = (~(Rbyx84 | Ittx84));
	assign Iayx84 = (Ybyx84 & Fcyx84);
	assign Fcyx84 = (~(W7ux84 | Mcyx84));
	assign Ybyx84 = (Tcyx84 & Adyx84);
	assign L8yx84 = (~(Hdyx84 & Uurx84));
	assign Hdyx84 = (F0wx84 & Odyx84);
	assign F0wx84 = (!Lwvx84);
	assign L1yx84 = (Vdyx84 & Me5w84);
	assign Vdyx84 = (Ceyx84 & Jeyx84);
	assign Jeyx84 = (~(Qeyx84 & Xeyx84));
	assign Xeyx84 = (~(Efyx84 & Uurx84));
	assign Uurx84 = (Zwvx84 & Lfyx84);
	assign Zwvx84 = (Sfyx84 | Zfyx84);
	assign Efyx84 = (~(Lwvx84 | Ggyx84));
	assign Ggyx84 = (!Uxvx84);
	assign Uxvx84 = (Fgux84 | Zfyx84);
	assign Lwvx84 = (Ngyx84 & Ugyx84);
	assign Qeyx84 = (~(Bhyx84 & Ihyx84));
	assign Ihyx84 = (Phyx84 & D8ux84);
	assign Phyx84 = (~(Znxx84 | Rqxx84));
	assign Znxx84 = (!Suxx84);
	assign Bhyx84 = (Whyx84 & Diyx84);
	assign Whyx84 = (F5yx84 ? Riyx84 : Kiyx84);
	assign Riyx84 = (Yiyx84 & Fjyx84);
	assign Fjyx84 = (~(W7ux84 | Mjyx84));
	assign Yiyx84 = (Tjyx84 & Adyx84);
	assign Kiyx84 = (Akyx84 & Hkyx84);
	assign Hkyx84 = (Okyx84 & Vkyx84);
	assign Akyx84 = (~(Clyx84 | Jlyx84));
	assign Ceyx84 = (~(Qlyx84 & Xlyx84));
	assign Qlyx84 = (~(Emyx84 & Lmyx84));
	assign Lmyx84 = (Smyx84 & Zmyx84);
	assign Zmyx84 = (~(Uvxx84 | Gnyx84));
	assign Smyx84 = (~(Nnyx84 | Unyx84));
	assign Emyx84 = (Boyx84 & Ioyx84);
	assign Ioyx84 = (~(Poyx84 | C4ux84));
	assign C4ux84 = (Kpyx84 ? Dpyx84 : Woyx84);
	assign Kpyx84 = (Rpyx84 & Ypyx84);
	assign Ypyx84 = (~(Fqyx84 & Mqyx84));
	assign Mqyx84 = (Tqyx84 | Aryx84);
	assign Rpyx84 = (Hryx84 | Aryx84);
	assign Dpyx84 = (F5yx84 ? Jlyx84 : Oryx84);
	assign Boyx84 = (Vryx84 & Csyx84);
	assign X0yx84 = (~(Jsyx84 & Qsyx84));
	assign Qsyx84 = (Xsyx84 & Etyx84);
	assign Etyx84 = (Ltyx84 & Styx84);
	assign Styx84 = (Ztyx84 & Guyx84);
	assign Guyx84 = (Nuyx84 & Xlrx84);
	assign Xlrx84 = (~(Uuyx84 & Bvyx84));
	assign Uuyx84 = (Si63a4 ? Pvyx84 : Ivyx84);
	assign Nuyx84 = (Rbrx84 & Kosx84);
	assign Kosx84 = (~(Wvyx84 & Dwyx84));
	assign Wvyx84 = (Ag63a4 ? Pvyx84 : Ivyx84);
	assign Rbrx84 = (~(Kwyx84 & Rwyx84));
	assign Kwyx84 = (Ei63a4 ? Pvyx84 : Ivyx84);
	assign Ztyx84 = (N2rx84 & Pwqx84);
	assign Pwqx84 = (~(Ywyx84 & Fxyx84));
	assign Ywyx84 = (Xh63a4 ? Pvyx84 : Ivyx84);
	assign N2rx84 = (~(Mxyx84 & Txyx84));
	assign Mxyx84 = (Zi63a4 ? Pvyx84 : Ivyx84);
	assign Ltyx84 = (Ayyx84 & Hyyx84);
	assign Hyyx84 = (F3tx84 & Ihrx84);
	assign Ihrx84 = (~(Oyyx84 & Vyyx84));
	assign Oyyx84 = (Li63a4 ? Pvyx84 : Ivyx84);
	assign F3tx84 = (~(Czyx84 & Jzyx84));
	assign Czyx84 = (Hg63a4 ? Pvyx84 : Ivyx84);
	assign Ayyx84 = (Vjsx84 & Nfsx84);
	assign Nfsx84 = (~(Qzyx84 & Xzyx84));
	assign Qzyx84 = (Jh63a4 ? Pvyx84 : Ivyx84);
	assign Vjsx84 = (~(E0zx84 & L0zx84));
	assign E0zx84 = (Qh63a4 ? Pvyx84 : Ivyx84);
	assign Xsyx84 = (S0zx84 & Z0zx84);
	assign Z0zx84 = (G1zx84 & N1zx84);
	assign N1zx84 = (U1zx84 & Yasx84);
	assign Yasx84 = (~(B2zx84 & I2zx84));
	assign B2zx84 = (Vg63a4 ? Pvyx84 : Ivyx84);
	assign U1zx84 = (Ieux84 & Wusx84);
	assign Wusx84 = (~(P2zx84 & W2zx84));
	assign P2zx84 = (O87w84 ? Pvyx84 : Ivyx84);
	assign Ieux84 = (~(D3zx84 & K3zx84));
	assign D3zx84 = (Ch63a4 ? Pvyx84 : Ivyx84);
	assign G1zx84 = (R3zx84 & C6sx84);
	assign C6sx84 = (~(Y3zx84 & F4zx84));
	assign Y3zx84 = (Og63a4 ? Pvyx84 : Ivyx84);
	assign R3zx84 = (~(Rdpx84 & M4zx84));
	assign M4zx84 = (~(T4zx84 & A5zx84));
	assign A5zx84 = (H5zx84 & O5zx84);
	assign O5zx84 = (V5zx84 & C6zx84);
	assign C6zx84 = (~(J6zx84 | Qp63a4[2]));
	assign J6zx84 = (Qp63a4[3] | Qp63a4[7]);
	assign V5zx84 = (~(Qp63a4[27] | Qp63a4[28]));
	assign H5zx84 = (Q6zx84 & X6zx84);
	assign X6zx84 = (~(Qp63a4[25] | Qp63a4[26]));
	assign Q6zx84 = (~(Qp63a4[22] | Qp63a4[23]));
	assign T4zx84 = (E7zx84 & L7zx84);
	assign L7zx84 = (S7zx84 & Z7zx84);
	assign Z7zx84 = (~(G8zx84 | Qp63a4[16]));
	assign G8zx84 = (Qp63a4[20] | Qp63a4[21]);
	assign S7zx84 = (~(Qp63a4[14] | Qp63a4[15]));
	assign E7zx84 = (N8zx84 & U8zx84);
	assign U8zx84 = (~(Qp63a4[11] | Qp63a4[13]));
	assign N8zx84 = (~(Qp63a4[0] | Qp63a4[10]));
	assign S0zx84 = (B9zx84 & I9zx84);
	assign I9zx84 = (P9zx84 & W9zx84);
	assign W9zx84 = (~(Jmqx84 & Dazx84));
	assign Jmqx84 = (Gj63a4 ? Pvyx84 : Ivyx84);
	assign P9zx84 = (~(Sdtx84 & Kazx84));
	assign Kazx84 = (~(Razx84 & Yazx84));
	assign Yazx84 = (Fbzx84 & Mbzx84);
	assign Mbzx84 = (Tbzx84 & Aczx84);
	assign Aczx84 = (Hczx84 & E6tx84);
	assign Hczx84 = (~(Oczx84 | Vczx84));
	assign Tbzx84 = (~(Cdzx84 | W8tx84));
	assign Fbzx84 = (Jdzx84 & Qdzx84);
	assign Qdzx84 = (~(Xdzx84 | Eezx84));
	assign Jdzx84 = (~(Lezx84 | Sezx84));
	assign Razx84 = (Zezx84 & Gfzx84);
	assign Gfzx84 = (Nfzx84 & Ufzx84);
	assign Ufzx84 = (~(Bgzx84 | Igzx84));
	assign Nfzx84 = (~(Pgzx84 | Wgzx84));
	assign Zezx84 = (Dhzx84 & Khzx84);
	assign Khzx84 = (~(Rhzx84 | Yhzx84));
	assign Dhzx84 = (~(Fizx84 | Mizx84));
	assign B9zx84 = (Zdtx84 & Tizx84);
	assign Tizx84 = (Iusx84 | Ajzx84);
	assign Ajzx84 = (Hjzx84 & Ojzx84);
	assign Ojzx84 = (Vjzx84 & Ckzx84);
	assign Ckzx84 = (Jkzx84 & Qkzx84);
	assign Qkzx84 = (Xkzx84 & Elzx84);
	assign Elzx84 = (~(Ftax84 & Gj63a4));
	assign Gj63a4 = (~(Llzx84 ^ Slzx84));
	assign Llzx84 = (~(Zlzx84 & Gmzx84));
	assign Gmzx84 = (Nmzx84 & Umzx84);
	assign Umzx84 = (~(Tt6w84 & Bnzx84));
	assign Nmzx84 = (~(Inzx84 & Pq6w84));
	assign Zlzx84 = (Pnzx84 & Wnzx84);
	assign Wnzx84 = (~(Dozx84 & O16w84));
	assign Pnzx84 = (Kozx84 | Piqx84);
	assign Xkzx84 = (~(V1bx84 & Zi63a4));
	assign Zi63a4 = (~(Rozx84 ^ Slzx84));
	assign Rozx84 = (~(Yozx84 & Fpzx84));
	assign Fpzx84 = (H6rx84 | Kozx84);
	assign Yozx84 = (Mpzx84 & Tpzx84);
	assign Mpzx84 = (~(I86w84 & Dozx84));
	assign Jkzx84 = (Aqzx84 & Hqzx84);
	assign Hqzx84 = (~(T0bx84 & Si63a4));
	assign Si63a4 = (~(Oqzx84 ^ Slzx84));
	assign Oqzx84 = (~(Vqzx84 & Crzx84));
	assign Crzx84 = (Kozx84 | Ltrx84);
	assign Vqzx84 = (Jrzx84 & Tpzx84);
	assign Jrzx84 = (~(Ap6w84 & Dozx84));
	assign Aqzx84 = (~(A1bx84 & Li63a4));
	assign Li63a4 = (~(Qrzx84 ^ Slzx84));
	assign Qrzx84 = (~(Xrzx84 & Eszx84));
	assign Eszx84 = (Akrx84 | Kozx84);
	assign Xrzx84 = (Lszx84 & Tpzx84);
	assign Lszx84 = (~(Ln6w84 & Dozx84));
	assign Vjzx84 = (Sszx84 & Zszx84);
	assign Zszx84 = (Gtzx84 & Ntzx84);
	assign Ntzx84 = (~(H1bx84 & Ei63a4));
	assign Ei63a4 = (~(Utzx84 ^ Slzx84));
	assign Utzx84 = (~(Buzx84 & Iuzx84));
	assign Iuzx84 = (Lfrx84 | Kozx84);
	assign Buzx84 = (Puzx84 & Tpzx84);
	assign Puzx84 = (~(Wl6w84 & Dozx84));
	assign Gtzx84 = (~(C2bx84 & Xh63a4));
	assign Xh63a4 = (~(Wuzx84 ^ Slzx84));
	assign Wuzx84 = (~(Dvzx84 & Kvzx84));
	assign Kvzx84 = (Yxqx84 | Kozx84);
	assign Dvzx84 = (Rvzx84 & Yvzx84);
	assign Yvzx84 = (~(Q66w84 & Dozx84));
	assign Rvzx84 = (Tmox84 | Fwzx84);
	assign Sszx84 = (Mwzx84 & Twzx84);
	assign Twzx84 = (~(Gxax84 & Hg63a4));
	assign Hg63a4 = (E6tx84 ? Hxzx84 : Axzx84);
	assign Mwzx84 = (~(Iyax84 & Qh63a4));
	assign Qh63a4 = (~(Oxzx84 ^ Slzx84));
	assign Oxzx84 = (~(Vxzx84 & Cyzx84));
	assign Cyzx84 = (Nd6w84 ? Qyzx84 : Jyzx84);
	assign Jyzx84 = (~(Dozx84 & T7px84));
	assign Vxzx84 = (Xyzx84 & Tpzx84);
	assign Xyzx84 = (Xksx84 | Kozx84);
	assign Hjzx84 = (Ezzx84 & Lzzx84);
	assign Lzzx84 = (Szzx84 & Zzzx84);
	assign Zzzx84 = (G00y84 & N00y84);
	assign N00y84 = (~(Uxax84 & Ag63a4));
	assign Ag63a4 = (Lssx84 ? Hxzx84 : Axzx84);
	assign G00y84 = (~(Pyax84 & Jh63a4));
	assign Jh63a4 = (~(U00y84 ^ Slzx84));
	assign U00y84 = (B10y84 | I10y84);
	assign I10y84 = (Ba6w84 ? W10y84 : P10y84);
	assign P10y84 = (Dozx84 & T7px84);
	assign B10y84 = (~(D20y84 & Tpzx84));
	assign D20y84 = (Fisx84 | Kozx84);
	assign Szzx84 = (K20y84 & R20y84);
	assign R20y84 = (~(M0bx84 & Ch63a4));
	assign Ch63a4 = (~(Y20y84 ^ Slzx84));
	assign Y20y84 = (~(F30y84 & M30y84));
	assign M30y84 = (Vhux84 | Kozx84);
	assign F30y84 = (T30y84 & Tpzx84);
	assign T30y84 = (~(Pq6w84 & Dozx84));
	assign K20y84 = (~(Wyax84 & Vg63a4));
	assign Vg63a4 = (~(A40y84 ^ Slzx84));
	assign A40y84 = (~(H40y84 & O40y84));
	assign O40y84 = (Qdsx84 | Kozx84);
	assign H40y84 = (V40y84 & Tpzx84);
	assign V40y84 = (~(My6w84 & Dozx84));
	assign Ezzx84 = (C50y84 & J50y84);
	assign J50y84 = (W2zx84 | Pusx84);
	assign Pusx84 = (!O87w84);
	assign O87w84 = (Q50y84 | X50y84);
	assign Q50y84 = (Vxsx84 ? L60y84 : E60y84);
	assign C50y84 = (S60y84 & Z60y84);
	assign Z60y84 = (~(Dzax84 & Og63a4));
	assign Og63a4 = (~(G70y84 ^ Slzx84));
	assign G70y84 = (~(N70y84 & U70y84));
	assign U70y84 = (B9sx84 | Kozx84);
	assign B9sx84 = (!Pgzx84);
	assign N70y84 = (B80y84 & Tpzx84);
	assign B80y84 = (~(Xw6w84 & Dozx84));
	assign S60y84 = (~(Lwax84 & Tf63a4));
	assign Zdtx84 = (I80y84 & P80y84);
	assign P80y84 = (V9ax84 ? D90y84 : W80y84);
	assign D90y84 = (R90y84 ? K90y84 : Iusx84);
	assign W80y84 = (Zwax84 | Y90y84);
	assign I80y84 = (Fa0y84 & Kdpx84);
	assign Fa0y84 = (~(Om5w84 & Ma0y84));
	assign Jsyx84 = (Ta0y84 & Ab0y84);
	assign Ab0y84 = (Hb0y84 & Ob0y84);
	assign Ob0y84 = (Vb0y84 & Cc0y84);
	assign Cc0y84 = (Jc0y84 & Fepx84);
	assign Fepx84 = (Qc0y84 & Xc0y84);
	assign Xc0y84 = (Ed0y84 & Ld0y84);
	assign Ld0y84 = (Shpx84 | Sd0y84);
	assign Ed0y84 = (Zd0y84 & Ge0y84);
	assign Ge0y84 = (~(Ne0y84 & Ue0y84));
	assign Ue0y84 = (~(D8gx84 | Bf0y84));
	assign Ne0y84 = (Yk5w84 & If0y84);
	assign Zd0y84 = (~(Qp63a4[1] & Rdpx84));
	assign Qc0y84 = (Pf0y84 & Wf0y84);
	assign Wf0y84 = (~(Dg0y84 & Nj63a4[1]));
	assign Pf0y84 = (T67w84 ? Rg0y84 : Kg0y84);
	assign T67w84 = (~(Yg0y84 ^ Slzx84));
	assign Yg0y84 = (~(Fh0y84 & Mh0y84));
	assign Mh0y84 = (Sd0y84 | Kozx84);
	assign Fh0y84 = (Th0y84 & Ai0y84);
	assign Ai0y84 = (~(Hk6w84 & Hi0y84));
	assign Th0y84 = (~(Kr5w84 & Dozx84));
	assign Rg0y84 = (Oi0y84 ? K90y84 : Iusx84);
	assign Kg0y84 = (Kzax84 | Y90y84);
	assign Jc0y84 = (Ydpx84 & Ompx84);
	assign Ompx84 = (Vi0y84 & Cj0y84);
	assign Cj0y84 = (~(Nj63a4[3] & Dg0y84));
	assign Vi0y84 = (Ys8x84 ? Qj0y84 : Jj0y84);
	assign Ys8x84 = (~(Xj0y84 ^ Slzx84));
	assign Xj0y84 = (~(Ek0y84 & Lk0y84));
	assign Lk0y84 = (Sk0y84 & Zk0y84);
	assign Zk0y84 = (Hanx84 | Gl0y84);
	assign Sk0y84 = (~(Ln6w84 & Bnzx84));
	assign Ek0y84 = (Nl0y84 & Ul0y84);
	assign Ul0y84 = (~(Uu5w84 & Dozx84));
	assign Nl0y84 = (Tlpx84 | Kozx84);
	assign Qj0y84 = (Bm0y84 ? K90y84 : Iusx84);
	assign Jj0y84 = (Huax84 | Y90y84);
	assign Ydpx84 = (Im0y84 & Pm0y84);
	assign Pm0y84 = (Wm0y84 & Dn0y84);
	assign Dn0y84 = (~(Kn0y84 & Rn0y84));
	assign Rn0y84 = (~(D8gx84 | Wl6w84));
	assign Kn0y84 = (Nr4w84 & If0y84);
	assign Wm0y84 = (Shpx84 | Yn0y84);
	assign Im0y84 = (Fo0y84 & Mo0y84);
	assign Mo0y84 = (~(Dg0y84 & Nj63a4[0]));
	assign Fo0y84 = (Y47w84 ? Ap0y84 : To0y84);
	assign Y47w84 = (~(Hp0y84 ^ Slzx84));
	assign Hp0y84 = (~(Op0y84 & Vp0y84));
	assign Vp0y84 = (~(Si6w84 & Hi0y84));
	assign Op0y84 = (Yn0y84 | Kozx84);
	assign Ap0y84 = (Cq0y84 ? K90y84 : Iusx84);
	assign To0y84 = (J2bx84 | Y90y84);
	assign Vb0y84 = (F4sx84 & U1sx84);
	assign U1sx84 = (Jq0y84 & Qq0y84);
	assign Qq0y84 = (Xq0y84 & Kdpx84);
	assign Xq0y84 = (~(Qp63a4[18] & Rdpx84));
	assign Jq0y84 = (Er0y84 & Lr0y84);
	assign Lr0y84 = (Shpx84 | Sr0y84);
	assign Er0y84 = (Xaax84 ? Gs0y84 : Zr0y84);
	assign Gs0y84 = (Ns0y84 ? K90y84 : Iusx84);
	assign Zr0y84 = (Yzax84 | Y90y84);
	assign F4sx84 = (Us0y84 & Bt0y84);
	assign Bt0y84 = (It0y84 & Kdpx84);
	assign It0y84 = (~(Qp63a4[19] & Rdpx84));
	assign Us0y84 = (Pt0y84 & Wt0y84);
	assign Wt0y84 = (Shpx84 | Du0y84);
	assign Pt0y84 = (Qaax84 ? Ru0y84 : Ku0y84);
	assign Ru0y84 = (Yu0y84 ? K90y84 : Iusx84);
	assign Ku0y84 = (Rzax84 | Y90y84);
	assign Hb0y84 = (Fv0y84 & Mv0y84);
	assign Mv0y84 = (U9rx84 & Nipx84);
	assign Nipx84 = (Tv0y84 & Aw0y84);
	assign Aw0y84 = (Hw0y84 & Ow0y84);
	assign Ow0y84 = (Shpx84 | Vw0y84);
	assign Hw0y84 = (Cx0y84 & Kdpx84);
	assign Cx0y84 = (~(Qp63a4[5] & Rdpx84));
	assign Tv0y84 = (Jx0y84 & Qx0y84);
	assign Qx0y84 = (~(Nj63a4[5] & Dg0y84));
	assign Jx0y84 = (F8ax84 ? Ey0y84 : Xx0y84);
	assign Ey0y84 = (Ly0y84 ? K90y84 : Iusx84);
	assign Xx0y84 = (Ttax84 | Y90y84);
	assign U9rx84 = (Sy0y84 & Zy0y84);
	assign Zy0y84 = (Gz0y84 & Kdpx84);
	assign Gz0y84 = (~(Qp63a4[12] & Rdpx84));
	assign Sy0y84 = (Nz0y84 & Uz0y84);
	assign Uz0y84 = (Shpx84 | B01y84);
	assign Nz0y84 = (Jaax84 ? P01y84 : I01y84);
	assign P01y84 = (W01y84 ? K90y84 : Iusx84);
	assign I01y84 = (O1bx84 | Y90y84);
	assign Fv0y84 = (Ixpx84 & Frqx84);
	assign Frqx84 = (D11y84 & K11y84);
	assign K11y84 = (R11y84 & Kdpx84);
	assign R11y84 = (~(Qp63a4[8] & Rdpx84));
	assign D11y84 = (Y11y84 & F21y84);
	assign F21y84 = (Shpx84 | M21y84);
	assign Y11y84 = (T8ax84 ? A31y84 : T21y84);
	assign A31y84 = (H31y84 ? K90y84 : Iusx84);
	assign T21y84 = (Ysax84 | Y90y84);
	assign Ixpx84 = (O31y84 & V31y84);
	assign V31y84 = (C41y84 & Kdpx84);
	assign C41y84 = (~(Qp63a4[6] & Rdpx84));
	assign O31y84 = (J41y84 & Q41y84);
	assign Q41y84 = (Shpx84 | X41y84);
	assign J41y84 = (M8ax84 ? L51y84 : E51y84);
	assign L51y84 = (Mtax84 ? Iusx84 : K90y84);
	assign E51y84 = (Mtax84 | Y90y84);
	assign Ta0y84 = (S51y84 & Z51y84);
	assign Z51y84 = (G61y84 & N61y84);
	assign N61y84 = (Trqx84 & Gaqx84);
	assign Gaqx84 = (U61y84 & B71y84);
	assign B71y84 = (I71y84 & P71y84);
	assign P71y84 = (Shpx84 | W71y84);
	assign I71y84 = (D81y84 & Kdpx84);
	assign D81y84 = (~(Qp63a4[4] & Rdpx84));
	assign U61y84 = (K81y84 & R81y84);
	assign R81y84 = (~(Dg0y84 & Nj63a4[4]));
	assign K81y84 = (Y7ax84 ? F91y84 : Y81y84);
	assign F91y84 = (M91y84 ? K90y84 : Iusx84);
	assign Y81y84 = (Auax84 | Y90y84);
	assign Trqx84 = (T91y84 & Aa1y84);
	assign Aa1y84 = (Ha1y84 & Kdpx84);
	assign Ha1y84 = (~(Qp63a4[9] & Rdpx84));
	assign T91y84 = (Oa1y84 & Va1y84);
	assign Va1y84 = (Shpx84 | Cb1y84);
	assign Oa1y84 = (R7ax84 ? Qb1y84 : Jb1y84);
	assign Qb1y84 = (Xb1y84 ? K90y84 : Iusx84);
	assign Jb1y84 = (Rsax84 | Y90y84);
	assign G61y84 = (Tmvx84 & Jzrx84);
	assign Jzrx84 = (Ec1y84 & Lc1y84);
	assign Lc1y84 = (Sc1y84 & Kdpx84);
	assign Sc1y84 = (~(Qp63a4[17] & Rdpx84));
	assign Ec1y84 = (Zc1y84 & Gd1y84);
	assign Gd1y84 = (Shpx84 | Nd1y84);
	assign Zc1y84 = (Caax84 ? Be1y84 : Ud1y84);
	assign Be1y84 = (Ie1y84 ? K90y84 : Iusx84);
	assign Ud1y84 = (F0bx84 | Y90y84);
	assign Tmvx84 = (Pe1y84 & We1y84);
	assign We1y84 = (Df1y84 & Kdpx84);
	assign Df1y84 = (~(Qp63a4[24] & Rdpx84));
	assign Pe1y84 = (Kf1y84 & Rf1y84);
	assign Rf1y84 = (Shpx84 | Yf1y84);
	assign Shpx84 = (!Sdtx84);
	assign Kf1y84 = (O9ax84 ? Mg1y84 : Fg1y84);
	assign Mg1y84 = (Tg1y84 ? K90y84 : Iusx84);
	assign Fg1y84 = (Byax84 | Y90y84);
	assign S51y84 = (Ah1y84 & Hh1y84);
	assign Hh1y84 = (Bmtx84 & Fotx84);
	assign Fotx84 = (Oh1y84 & Vh1y84);
	assign Vh1y84 = (Ci1y84 & Ji1y84);
	assign Ji1y84 = (~(Eo5w84 & Ma0y84));
	assign Ci1y84 = (Qi1y84 & Kdpx84);
	assign Qi1y84 = (~(Qp63a4[30] & Rdpx84));
	assign Oh1y84 = (Xi1y84 & Ej1y84);
	assign Ej1y84 = (~(Sdtx84 & Dwdx84));
	assign Xi1y84 = (H9ax84 ? Sj1y84 : Lj1y84);
	assign Sj1y84 = (Zj1y84 ? K90y84 : Iusx84);
	assign Lj1y84 = (Ouax84 | Y90y84);
	assign Bmtx84 = (Gk1y84 & Nk1y84);
	assign Nk1y84 = (Uk1y84 & Bl1y84);
	assign Bl1y84 = (~(Ma0y84 & Th5w84));
	assign Uk1y84 = (Il1y84 & Kdpx84);
	assign Il1y84 = (~(Qp63a4[29] & Rdpx84));
	assign Gk1y84 = (Pl1y84 & Wl1y84);
	assign Wl1y84 = (~(Sdtx84 & Vitx84));
	assign Pl1y84 = (A9ax84 ? Km1y84 : Dm1y84);
	assign Km1y84 = (Rm1y84 ? K90y84 : Iusx84);
	assign Dm1y84 = (Swax84 | Y90y84);
	assign Ah1y84 = (H0xx84 & Ehpx84);
	assign Ehpx84 = (Ym1y84 & Fn1y84);
	assign Fn1y84 = (~(Nj63a4[2] & Dg0y84));
	assign Dg0y84 = (Mn1y84 & If0y84);
	assign Mn1y84 = (~(Tn1y84 | Ap6w84));
	assign Ym1y84 = (Ao1y84 & Ho1y84);
	assign Ho1y84 = (~(Oo1y84 & Vo1y84));
	assign Vo1y84 = (~(Ambx84 | Ewax84));
	assign Oo1y84 = (Hj5w84 & I5bx84);
	assign Ao1y84 = (~(Cp1y84 & Ascx84));
	assign Cp1y84 = (Tf63a4 ? Pvyx84 : Ivyx84);
	assign Tf63a4 = (~(Jp1y84 ^ Slzx84));
	assign Jp1y84 = (~(Qp1y84 & Xp1y84));
	assign Xp1y84 = (Eq1y84 & Lq1y84);
	assign Lq1y84 = (~(Wl6w84 & Hi0y84));
	assign Hi0y84 = (Sq1y84 | Bnzx84);
	assign Sq1y84 = (~(Zq1y84 & Gr1y84));
	assign Gr1y84 = (~(Nr1y84 & Ur1y84));
	assign Ur1y84 = (~(Wbcx84 | Pqbx84));
	assign Nr1y84 = (~(Bs1y84 | Xvax84));
	assign Zq1y84 = (~(Is1y84 & I5bx84));
	assign Is1y84 = (~(G4bx84 | Evix84));
	assign Eq1y84 = (Tn1y84 | Gl0y84);
	assign Qp1y84 = (Ps1y84 & Ws1y84);
	assign Ws1y84 = (~(Ct5w84 & Dozx84));
	assign Ps1y84 = (Zhpx84 | Kozx84);
	assign H0xx84 = (~(Aaux84 | Me5w84));
	assign Aaux84 = (~(Dt1y84 & Kt1y84));
	assign Kt1y84 = (Rt1y84 & Yt1y84);
	assign Yt1y84 = (~(Up5w84 & Ma0y84));
	assign Ma0y84 = (Auvx84 & If0y84);
	assign If0y84 = (Fu1y84 & Ol2x84);
	assign Fu1y84 = (J0dx84 & Ambx84);
	assign Auvx84 = (~(Wl6w84 | Ap6w84));
	assign Rt1y84 = (Mu1y84 & Kdpx84);
	assign Kdpx84 = (~(Tu1y84 & Ol2x84));
	assign Mu1y84 = (~(Qp63a4[31] & Rdpx84));
	assign Rdpx84 = (~(Av1y84 & Hv1y84));
	assign Hv1y84 = (~(Ol2x84 & Ov1y84));
	assign Ov1y84 = (Vv1y84 | Cw1y84);
	assign Cw1y84 = (Tq2x84 ? Gz4w84 : Jw1y84);
	assign Jw1y84 = (~(Qw1y84 | D4dx84));
	assign Vv1y84 = (~(Xw1y84 & Ex1y84));
	assign Ex1y84 = (~(Lx1y84 & Ambx84));
	assign Lx1y84 = (~(Sx1y84 & Zx1y84));
	assign Zx1y84 = (Fn2x84 | Ns2x84);
	assign Sx1y84 = (Gy1y84 & Naxx84);
	assign Gy1y84 = (Ny1y84 | Uy1y84);
	assign Av1y84 = (Bz1y84 & Iz1y84);
	assign Bz1y84 = (~(I5bx84 & Pz1y84));
	assign Pz1y84 = (~(Wz1y84 & D02y84));
	assign D02y84 = (Yshx84 | Ewax84);
	assign Wz1y84 = (Qxmx84 | Evix84);
	assign Dt1y84 = (K02y84 & R02y84);
	assign R02y84 = (~(Sdtx84 & Ysvx84));
	assign Sdtx84 = (Y02y84 & Ol2x84);
	assign Y02y84 = (~(Fmvx84 | Kzvx84));
	assign K02y84 = (Gqax84 ? M12y84 : F12y84);
	assign M12y84 = (O7xx84 ? K90y84 : Iusx84);
	assign K90y84 = (!Pvyx84);
	assign Pvyx84 = (~(T12y84 & A22y84));
	assign A22y84 = (H22y84 & O22y84);
	assign T12y84 = (V22y84 & C32y84);
	assign C32y84 = (~(I5bx84 & Y6bx84));
	assign V22y84 = (P1mx84 | Zo2x84);
	assign F12y84 = (J32y84 | Y90y84);
	assign Y90y84 = (!Ivyx84);
	assign Ivyx84 = (~(Q32y84 & H22y84));
	assign H22y84 = (~(Ol2x84 & X32y84));
	assign X32y84 = (~(E42y84 & L42y84));
	assign E42y84 = (S42y84 & Z42y84);
	assign Z42y84 = (~(G52y84 & N52y84));
	assign N52y84 = (N4ix84 | C0dx84);
	assign S42y84 = (~(Hwmx84 & Ambx84));
	assign Q32y84 = (Iusx84 & O22y84);
	assign Iusx84 = (~(U52y84 & Devx84));
	assign U52y84 = (I5bx84 & Ambx84);
	assign Pwxx84 = (~(Tlwx84 | Q66w84));
	assign Kywx84 = (B62y84 & Leex84);
	assign B62y84 = (~(L4ox84 & I62y84));
	assign I62y84 = (J8cx84 | Fcdx84);
	assign Wxwx84 = (~(C2ix84 & P62y84));
	assign P62y84 = (~(W62y84 & D72y84));
	assign D72y84 = (~(K72y84 | E9cx84));
	assign K72y84 = (R72y84 & Y72y84);
	assign Y72y84 = (F82y84 & Qklx84);
	assign F82y84 = (~(Ey5w84 | Wz5w84));
	assign R72y84 = (M82y84 & Ihdx84);
	assign M82y84 = (T82y84 & I86w84);
	assign W62y84 = (Nd6w84 & A92y84);
	assign A92y84 = (Ifmx84 | Q66w84);
	assign Vtwx84 = (H92y84 & O92y84);
	assign O92y84 = (~(V92y84 & Uj2x84));
	assign V92y84 = (~(Jxmx84 | B3dx84));
	assign H92y84 = (~(Ca2y84 & Qxmx84));
	assign Ca2y84 = (~(Ja2y84 & Qa2y84));
	assign Qa2y84 = (Xa2y84 & Eb2y84);
	assign Eb2y84 = (~(Lb2y84 & A2ox84));
	assign Xa2y84 = (J9bx84 | Hgvx84);
	assign Ja2y84 = (~(Sb2y84 | Zb2y84));
	assign Zb2y84 = (~(Y4dx84 | Wbcx84));
	assign Sb2y84 = (Yqcx84 ? Nc2y84 : Gc2y84);
	assign Nc2y84 = (Eelx84 & Rvlx84);
	assign Wqwx84 = (Uc2y84 & Bd2y84);
	assign Bd2y84 = (Id2y84 & Urnx84);
	assign Urnx84 = (Pd2y84 & Wd2y84);
	assign Wd2y84 = (Gqox84 | Ambx84);
	assign Id2y84 = (De2y84 & Mi42a4);
	assign Mi42a4 = (~(Ti42a4 & H6dx84));
	assign Ti42a4 = (~(Aj42a4 & Hj42a4));
	assign Hj42a4 = (Oj42a4 & Vj42a4);
	assign Vj42a4 = (~(Xgwx84 & Ck42a4));
	assign Ck42a4 = (~(Jk42a4 & Qk42a4));
	assign Qk42a4 = (~(Xk42a4 & El42a4));
	assign Xk42a4 = (~(M6xx84 | Wqbx84));
	assign Jk42a4 = (Bqwx84 | Hu2x84);
	assign Oj42a4 = (~(Gf6w84 & Ll42a4));
	assign Ll42a4 = (~(Sl42a4 & Zl42a4));
	assign Zl42a4 = (~(Gm42a4 & Nm42a4));
	assign Nm42a4 = (Lzlx84 & Um42a4);
	assign Gm42a4 = (Momx84 & Bn42a4);
	assign Sl42a4 = (!Ejnx84);
	assign Aj42a4 = (In42a4 & Pn42a4);
	assign Pn42a4 = (~(L2cx84 & Wn42a4));
	assign In42a4 = (~(Pxbx84 & Do42a4));
	assign Do42a4 = (~(Ko42a4 & Ro42a4));
	assign Ro42a4 = (Yo42a4 & Fp42a4);
	assign Fp42a4 = (Mp42a4 | M6xx84);
	assign Mp42a4 = (!Tp42a4);
	assign Yo42a4 = (~(Nzfx84 | Aq42a4));
	assign Nzfx84 = (Hq42a4 & W05w84);
	assign Hq42a4 = (~(M6xx84 | Gf6w84));
	assign Ko42a4 = (Oq42a4 & Vq42a4);
	assign Vq42a4 = (~(Uacx84 & Devx84));
	assign Oq42a4 = (~(Nacx84 & E3wx84));
	assign De2y84 = (~(Dzox84 & Pxbx84));
	assign Uc2y84 = (~(Cr42a4 | Jr42a4));
	assign Cr42a4 = (Bw2x84 ? Rfnx84 : Ljnx84);
	assign Ljnx84 = (Qr42a4 & Iqbx84);
	assign Qr42a4 = (~(Ambx84 | G4wx84));
	assign Cf4x84 = (~(Xr42a4 & Es42a4));
	assign Es42a4 = (~(HREADY & Ls42a4));
	assign Ls42a4 = (~(Ss42a4 & Zs42a4));
	assign Zs42a4 = (Gt42a4 & Nt42a4);
	assign Nt42a4 = (Ut42a4 & Bu42a4);
	assign Bu42a4 = (Iu42a4 & P5wx84);
	assign Ut42a4 = (Pu42a4 & Wu42a4);
	assign Wu42a4 = (~(Dv42a4 & Kv42a4));
	assign Kv42a4 = (Plnx84 & Ns2x84);
	assign Dv42a4 = (~(Rv42a4 | Yv42a4));
	assign Pu42a4 = (~(Fw42a4 & W05w84));
	assign Fw42a4 = (Zg6w84 & Mw42a4);
	assign Mw42a4 = (~(Tw42a4 & Ax42a4));
	assign Ax42a4 = (~(Ilnx84 & Pxbx84));
	assign Tw42a4 = (~(Hx42a4 | Atix84));
	assign Gt42a4 = (Ox42a4 & Vx42a4);
	assign Vx42a4 = (Cy42a4 & Jy42a4);
	assign Jy42a4 = (~(Qy42a4 & Cavx84));
	assign Qy42a4 = (~(Raex84 | Hgvx84));
	assign Cy42a4 = (~(Xy42a4 & Ffox84));
	assign Xy42a4 = (~(Yxcx84 | Hu2x84));
	assign Ox42a4 = (Ez42a4 & Lz42a4);
	assign Lz42a4 = (~(Sz42a4 & Zz42a4));
	assign Zz42a4 = (~(U4wx84 & G052a4));
	assign G052a4 = (Jxmx84 | N052a4);
	assign U4wx84 = (!U052a4);
	assign Ez42a4 = (~(U8lx84 & B152a4));
	assign B152a4 = (~(V9ox84 & I152a4));
	assign I152a4 = (Yxcx84 | Nbix84);
	assign Yxcx84 = (!Eelx84);
	assign Ss42a4 = (P152a4 & W152a4);
	assign W152a4 = (D252a4 & K252a4);
	assign K252a4 = (R252a4 & Y252a4);
	assign Y252a4 = (~(Gc2y84 & F352a4));
	assign R252a4 = (~(Ilnx84 & Xgwx84));
	assign Ilnx84 = (~(M6xx84 | P1mx84));
	assign D252a4 = (M352a4 & T352a4);
	assign T352a4 = (~(A452a4 & H6dx84));
	assign A452a4 = (~(H452a4 & O452a4));
	assign O452a4 = (V452a4 & C552a4);
	assign C552a4 = (~(C2ix84 & J552a4));
	assign J552a4 = (~(Q552a4 & X552a4));
	assign X552a4 = (~(Jpnx84 & Ub6w84));
	assign Q552a4 = (E652a4 & L652a4);
	assign L652a4 = (~(S652a4 & Z652a4));
	assign Z652a4 = (G752a4 & X8cx84);
	assign G752a4 = (~(Wcbx84 | Y46w84));
	assign S652a4 = (Momx84 & N752a4);
	assign E652a4 = (~(L6mx84 & U752a4));
	assign U752a4 = (~(B852a4 & I852a4));
	assign I852a4 = (P852a4 & W852a4);
	assign W852a4 = (~(D952a4 & Mcdx84));
	assign D952a4 = (~(Q1xx84 | Qzkx84));
	assign P852a4 = (~(K952a4 & Ubwx84));
	assign K952a4 = (~(R952a4 | Ba6w84));
	assign B852a4 = (Y952a4 & Fa52a4);
	assign Fa52a4 = (~(Nd6w84 & Ma52a4));
	assign Ma52a4 = (~(Ta52a4 & Ab52a4));
	assign Ab52a4 = (Q1cx84 | Hb52a4);
	assign Ta52a4 = (Ob52a4 & Vb52a4);
	assign Vb52a4 = (~(Cc52a4 & Zfdx84));
	assign Cc52a4 = (~(R952a4 | Ey5w84));
	assign Ob52a4 = (~(Jc52a4 & Ihdx84));
	assign Jc52a4 = (~(Bhdx84 | Iicx84));
	assign Y952a4 = (Y46w84 ? Xc52a4 : Qc52a4);
	assign Xc52a4 = (~(Tlwx84 & Wcbx84));
	assign Qc52a4 = (~(Lfdx84 & Gwbx84));
	assign V452a4 = (Ed52a4 & Ld52a4);
	assign Ld52a4 = (~(Sd52a4 & Huhx84));
	assign Sd52a4 = (~(Xlkx84 | J8cx84));
	assign Ed52a4 = (~(Zd52a4 & Aq42a4));
	assign Zd52a4 = (~(Fmvx84 | Yrbx84));
	assign H452a4 = (~(Ge52a4 | Ne52a4));
	assign Ne52a4 = (Hu2x84 ? Bf52a4 : Ue52a4);
	assign Ue52a4 = (~(Vkdx84 | Gz4w84));
	assign Vkdx84 = (!Jsrx84);
	assign Ge52a4 = (~(If52a4 & Pf52a4));
	assign Pf52a4 = (~(Wf52a4 & F3mx84));
	assign Wf52a4 = (~(Dg52a4 & Kg52a4));
	assign Kg52a4 = (~(X7dx84 & Rg52a4));
	assign Rg52a4 = (~(Yg52a4 & Fh52a4));
	assign Fh52a4 = (Mh52a4 & Th52a4);
	assign Th52a4 = (N3cx84 | Y46w84);
	assign Mh52a4 = (Ai52a4 | Efdx84);
	assign Yg52a4 = (Gf6w84 & Hi52a4);
	assign Hi52a4 = (B4cx84 | Hb52a4);
	assign Dg52a4 = (Oi52a4 & Vi52a4);
	assign Vi52a4 = (~(Cj52a4 & Jj52a4));
	assign Cj52a4 = (S6mx84 & J8cx84);
	assign Oi52a4 = (~(X8cx84 & Qj52a4));
	assign Qj52a4 = (~(Xj52a4 & Ek52a4));
	assign Ek52a4 = (~(J5mx84 & Ixwx84));
	assign Xj52a4 = (Lk52a4 & C5mx84);
	assign If52a4 = (~(Iqbx84 & Y1gx84));
	assign M352a4 = (~(Sk52a4 & Gpbx84));
	assign Sk52a4 = (~(Zk52a4 & Gl52a4));
	assign Gl52a4 = (Nl52a4 & Ul52a4);
	assign Ul52a4 = (~(Bm52a4 & Vzcx84));
	assign Bm52a4 = (~(Im52a4 & Pm52a4));
	assign Pm52a4 = (~(Xhvx84 & E3wx84));
	assign Im52a4 = (Hkdx84 | Bw2x84);
	assign Nl52a4 = (Wm52a4 & Dn52a4);
	assign Wm52a4 = (~(Kn52a4 & Nacx84));
	assign Kn52a4 = (~(S1dx84 | Qxmx84));
	assign Zk52a4 = (Rn52a4 & Yn52a4);
	assign Yn52a4 = (Qldx84 | Ewax84);
	assign Qldx84 = (!Fo52a4);
	assign Rn52a4 = (~(Mo52a4 & Pqbx84));
	assign Mo52a4 = (~(To52a4 & Ebox84));
	assign To52a4 = (~(Y6bx84 | Ap52a4));
	assign P152a4 = (Hp52a4 & Op52a4);
	assign Op52a4 = (Yrbx84 ? Cq52a4 : Vp52a4);
	assign Cq52a4 = (~(Ogvx84 & E3wx84));
	assign Vp52a4 = (~(Jq52a4 & Pxbx84));
	assign Hp52a4 = (~(Jr42a4 | Qq52a4));
	assign Qq52a4 = (Zvix84 & Rfnx84);
	assign Jr42a4 = (~(Cubx84 & Xq52a4));
	assign Xq52a4 = (J9bx84 | Jnix84);
	assign Xr42a4 = (Er52a4 & Lr52a4);
	assign Lr52a4 = (~(Sr52a4 & Qoox84));
	assign Sr52a4 = (~(O8bx84 | Evix84));
	assign Er52a4 = (~(Zo2x84 & Zr52a4));
	assign Zr52a4 = (Wpcx84 | Hbmx84);
	assign We4x84 = (Gs52a4 & Ns52a4);
	assign Ns52a4 = (~(Us52a4 & Bt52a4));
	assign Bt52a4 = (It52a4 & Pt52a4);
	assign Pt52a4 = (Wt52a4 & Du52a4);
	assign Du52a4 = (Ku52a4 & Ru52a4);
	assign Ku52a4 = (~(Yu52a4 & Fv52a4));
	assign Fv52a4 = (~(Xtcx84 | Nd6w84));
	assign Yu52a4 = (Mv52a4 & Q66w84);
	assign Wt52a4 = (Tv52a4 & Aw52a4);
	assign Aw52a4 = (~(Hw52a4 & Ow52a4));
	assign Ow52a4 = (~(Yshx84 | J13x84));
	assign Hw52a4 = (Mlbx84 & O1px84);
	assign Tv52a4 = (~(Vw52a4 & Huox84));
	assign Huox84 = (Cx52a4 & Xgwx84);
	assign Cx52a4 = (~(Qtcx84 | Vx2x84));
	assign Vw52a4 = (Hwmx84 & Rufx84);
	assign Rufx84 = (!Mw5w84);
	assign It52a4 = (Jx52a4 & Qx52a4);
	assign Qx52a4 = (~(Xhvx84 & Gwix84));
	assign Xhvx84 = (Zvix84 & H6dx84);
	assign Jx52a4 = (Xx52a4 & Ey52a4);
	assign Ey52a4 = (~(Ly52a4 & Phdx84));
	assign Ly52a4 = (~(B5bx84 | Tswx84));
	assign Xx52a4 = (~(Pz2x84 & Sy52a4));
	assign Sy52a4 = (~(Zy52a4 & Gz52a4));
	assign Gz52a4 = (~(Nz52a4 & Phdx84));
	assign Nz52a4 = (~(Mycx84 | N4bx84));
	assign Zy52a4 = (~(Zvix84 & Nwix84));
	assign Us52a4 = (Uz52a4 & B062a4);
	assign B062a4 = (I062a4 & P062a4);
	assign P062a4 = (~(W062a4 & H6dx84));
	assign W062a4 = (~(D162a4 & K162a4));
	assign K162a4 = (R162a4 & Y162a4);
	assign Y162a4 = (F262a4 & W3dx84);
	assign F262a4 = (~(M262a4 & Ovnx84));
	assign M262a4 = (T262a4 & A362a4);
	assign A362a4 = (~(Jmcx84 & H362a4));
	assign H362a4 = (~(O362a4 & Ai52a4));
	assign O362a4 = (G36w84 | Wz5w84);
	assign R162a4 = (V362a4 & C462a4);
	assign C462a4 = (~(Huhx84 & J462a4));
	assign J462a4 = (~(Q462a4 & X462a4));
	assign X462a4 = (~(E8dx84 & E562a4));
	assign E562a4 = (~(L562a4 & S562a4));
	assign S562a4 = (~(Z562a4 & Grnx84));
	assign Z562a4 = (~(Xlkx84 | O16w84));
	assign L562a4 = (~(G662a4 & Ihdx84));
	assign G662a4 = (Ixwx84 & S6mx84);
	assign Q462a4 = (L4ox84 | Ouhx84);
	assign V362a4 = (~(Yrbx84 & N662a4));
	assign N662a4 = (~(U662a4 & B762a4));
	assign B762a4 = (Ucox84 | Zbox84);
	assign Zbox84 = (Yqcx84 | Hu2x84);
	assign U662a4 = (~(Rzhx84 & Tsix84));
	assign D162a4 = (I762a4 & P762a4);
	assign P762a4 = (W762a4 & D862a4);
	assign D862a4 = (~(Ysox84 & Um42a4));
	assign Um42a4 = (Iicx84 ? Lfdx84 : N752a4);
	assign Ysox84 = (K862a4 & Grnx84);
	assign Grnx84 = (Bn42a4 & Gwbx84);
	assign K862a4 = (~(Mebx84 | Iokx84));
	assign Mebx84 = (~(F8ox84 & Edmx84));
	assign W762a4 = (Ucox84 | Evix84);
	assign I762a4 = (R862a4 & Y862a4);
	assign R862a4 = (Ba6w84 ? M962a4 : F962a4);
	assign M962a4 = (~(T962a4 & Y46w84));
	assign T962a4 = (Fcdx84 & Wadx84);
	assign F962a4 = (~(Mv52a4 & L2cx84));
	assign I062a4 = (Aa62a4 & Ha62a4);
	assign Ha62a4 = (~(Oa62a4 & Qxmx84));
	assign Oa62a4 = (~(Va62a4 & Cb62a4));
	assign Cb62a4 = (~(Ffox84 & Tsix84));
	assign Va62a4 = (Jb62a4 & V9ox84);
	assign V9ox84 = (!Cxfx84);
	assign Cxfx84 = (Teix84 & Wqbx84);
	assign Jb62a4 = (~(Qb62a4 & Mlbx84));
	assign Qb62a4 = (~(Rybx84 | Ewax84));
	assign Aa62a4 = (~(Xb62a4 & Hgvx84));
	assign Xb62a4 = (~(Ec62a4 & Lc62a4));
	assign Lc62a4 = (~(Sc62a4 & N052a4));
	assign Ec62a4 = (Zc62a4 & Gd62a4);
	assign Gd62a4 = (~(Nd62a4 & Gwix84));
	assign Nd62a4 = (~(Fycx84 | Bw2x84));
	assign Zc62a4 = (~(Tq2x84 & Ud62a4));
	assign Ud62a4 = (~(Be62a4 & Ie62a4));
	assign Ie62a4 = (~(Pe62a4 & M0px84));
	assign Pe62a4 = (~(Lrfx84 | Eelx84));
	assign Eelx84 = (~(We62a4 | Qq8x84));
	assign Be62a4 = (~(Zvix84 & J13x84));
	assign Uz52a4 = (Df62a4 & Kf62a4);
	assign Df62a4 = (Rf62a4 & Yf62a4);
	assign Yf62a4 = (~(Rzhx84 & O8px84));
	assign Rf62a4 = (Fg62a4 | Mg62a4);
	assign Gs52a4 = (Bw2x84 | HREADY);
	assign Qe4x84 = (Tg62a4 & Ah62a4);
	assign Ah62a4 = (~(Hh62a4 & Oh62a4));
	assign Oh62a4 = (Vh62a4 & Ci62a4);
	assign Ci62a4 = (Ji62a4 & Qi62a4);
	assign Qi62a4 = (Xi62a4 & Iu42a4);
	assign Xi62a4 = (Ru52a4 & Cubx84);
	assign Ru52a4 = (~(A7cx84 & J0dx84));
	assign Ji62a4 = (Ej62a4 & Lj62a4);
	assign Lj62a4 = (~(Sj62a4 & U052a4));
	assign U052a4 = (N4ix84 & G4bx84);
	assign Sj62a4 = (~(Yrix84 | Yrbx84));
	assign Ej62a4 = (~(Zj62a4 & X8cx84));
	assign Zj62a4 = (~(E2cx84 | Y46w84));
	assign Vh62a4 = (Gk62a4 & Nk62a4);
	assign Nk62a4 = (Uk62a4 & Bl62a4);
	assign Bl62a4 = (~(Momx84 & Il62a4));
	assign Il62a4 = (~(I4cx84 & Pl62a4));
	assign Pl62a4 = (~(Oxlx84 & Wl62a4));
	assign Wl62a4 = (~(Dm62a4 & Q66w84));
	assign Dm62a4 = (Km62a4 & Pxwx84);
	assign Pxwx84 = (!Lfdx84);
	assign Km62a4 = (Eobx84 | G36w84);
	assign Uk62a4 = (~(Undx84 & Rm62a4));
	assign Rm62a4 = (~(B0gx84 & Ym62a4));
	assign Ym62a4 = (Wtfx84 | H6dx84);
	assign Wtfx84 = (!Javx84);
	assign Javx84 = (Bw2x84 & G4bx84);
	assign Gk62a4 = (Fn62a4 & Mn62a4);
	assign Mn62a4 = (~(Tn62a4 & Y1gx84));
	assign Fn62a4 = (Ao62a4 | Ns2x84);
	assign Hh62a4 = (Ho62a4 & Oo62a4);
	assign Oo62a4 = (Vo62a4 & Cp62a4);
	assign Cp62a4 = (Jp62a4 & Qp62a4);
	assign Qp62a4 = (~(Xp62a4 & Gpbx84));
	assign Xp62a4 = (~(Eq62a4 & Lq62a4));
	assign Lq62a4 = (~(Sq62a4 & Vx2x84));
	assign Eq62a4 = (Zq62a4 & Gr62a4);
	assign Gr62a4 = (~(Tn62a4 & Nr62a4));
	assign Zq62a4 = (~(Hwmx84 & Ur62a4));
	assign Ur62a4 = (~(Bs62a4 & Plnx84));
	assign Bs62a4 = (~(W05w84 | Mw5w84));
	assign Jp62a4 = (Is62a4 & Ps62a4);
	assign Ps62a4 = (~(Ws62a4 & Dt62a4));
	assign Is62a4 = (~(X7dx84 & Kt62a4));
	assign Kt62a4 = (~(Rt62a4 & Yt62a4));
	assign Yt62a4 = (Wcbx84 | G36w84);
	assign Rt62a4 = (Fu62a4 & Hb52a4);
	assign Fu62a4 = (~(Mu62a4 & Z6mx84));
	assign Mu62a4 = (R952a4 | Y46w84);
	assign Vo62a4 = (Tu62a4 & Av62a4);
	assign Av62a4 = (~(Pxbx84 & Hv62a4));
	assign Hv62a4 = (~(Ov62a4 & Vv62a4));
	assign Vv62a4 = (~(Cw62a4 | F7bx84));
	assign Cw62a4 = (Jw62a4 & Yrbx84);
	assign Jw62a4 = (Qw62a4 & Ewax84);
	assign Qw62a4 = (F2gx84 | Xw62a4);
	assign Ov62a4 = (Ex62a4 & Lx62a4);
	assign Lx62a4 = (~(Fn2x84 & Sx62a4));
	assign Sx62a4 = (~(Ny1y84 & Zx62a4));
	assign Zx62a4 = (Wbcx84 | Pqbx84);
	assign Ex62a4 = (Zo2x84 ? Ny62a4 : Gy62a4);
	assign Ny62a4 = (Qxmx84 & Uy62a4);
	assign Uy62a4 = (Mmvx84 | Yybx84);
	assign Gy62a4 = (S1dx84 | Hu2x84);
	assign Tu62a4 = (~(Ykwx84 & Uacx84));
	assign Ho62a4 = (Bz62a4 & Iz62a4);
	assign Iz62a4 = (Dccx84 & Pz62a4);
	assign Pz62a4 = (Jxmx84 | P1mx84);
	assign Bz62a4 = (Wz62a4 & D072a4);
	assign Wz62a4 = (Gf6w84 ? R072a4 : K072a4);
	assign R072a4 = (Y072a4 & F172a4);
	assign F172a4 = (M172a4 | J8cx84);
	assign Y072a4 = (T172a4 & A272a4);
	assign A272a4 = (~(Gz4w84 & H272a4));
	assign H272a4 = (~(O272a4 & V272a4));
	assign V272a4 = (~(Oxlx84 & C372a4));
	assign C372a4 = (~(J372a4 & Y46w84));
	assign J372a4 = (~(Iicx84 | I86w84));
	assign O272a4 = (I4cx84 | Ixwx84);
	assign I4cx84 = (!X8cx84);
	assign T172a4 = (~(V1ix84 & Oxlx84));
	assign K072a4 = (Q372a4 & X372a4);
	assign X372a4 = (~(J5mx84 & E472a4));
	assign E472a4 = (Leex84 | Ba6w84);
	assign Q372a4 = (~(Ub6w84 & L472a4));
	assign L472a4 = (~(S472a4 & Z472a4));
	assign Z472a4 = (Z6mx84 | E2cx84);
	assign S472a4 = (~(G572a4 | J5mx84));
	assign G572a4 = (Momx84 & O16w84);
	assign Tg62a4 = (Vx2x84 | HREADY);
	assign Ke4x84 = (N572a4 & U572a4);
	assign U572a4 = (~(B672a4 & I672a4));
	assign I672a4 = (P672a4 & W672a4);
	assign W672a4 = (D772a4 & K772a4);
	assign K772a4 = (~(R772a4 & Sc62a4));
	assign R772a4 = (~(N052a4 | N4ix84));
	assign D772a4 = (A8ix84 & P5wx84);
	assign P5wx84 = (~(Rfnx84 & Gcvx84));
	assign P672a4 = (Y772a4 & F872a4);
	assign F872a4 = (~(M872a4 & Mlbx84));
	assign M872a4 = (Vx2x84 & T872a4);
	assign T872a4 = (Ozcx84 | Fo52a4);
	assign Y772a4 = (~(A972a4 & Rzhx84));
	assign A972a4 = (~(N4bx84 | Fn2x84));
	assign B672a4 = (H972a4 & O972a4);
	assign O972a4 = (V972a4 & Ca72a4);
	assign Ca72a4 = (~(Ja72a4 & Phdx84));
	assign V972a4 = (Qa72a4 & Xa72a4);
	assign Xa72a4 = (~(Eb72a4 & Gwix84));
	assign Eb72a4 = (~(H8px84 | Tsix84));
	assign Qa72a4 = (~(Kprx84 & Lb72a4));
	assign Lb72a4 = (~(Sb72a4 & Zb72a4));
	assign Zb72a4 = (~(Ogvx84 & U8lx84));
	assign Ogvx84 = (Gc72a4 & Tsix84);
	assign Sb72a4 = (~(Rzhx84 & O1px84));
	assign H972a4 = (Kf62a4 & Nc72a4);
	assign Nc72a4 = (~(Uc72a4 & H6dx84));
	assign Uc72a4 = (~(Bd72a4 & Id72a4));
	assign Id72a4 = (Pd72a4 & Wd72a4);
	assign Pd72a4 = (~(De72a4 & Ke72a4));
	assign Ke72a4 = (E8dx84 & Re72a4);
	assign Re72a4 = (~(Ye72a4 & Ff72a4));
	assign Ye72a4 = (Eobx84 ? Qzkx84 : Ai52a4);
	assign De72a4 = (X7dx84 & Ixwx84);
	assign Bd72a4 = (Y862a4 & Mf72a4);
	assign Y862a4 = (Tf72a4 & Ag72a4);
	assign Ag72a4 = (~(Hg72a4 & Ovnx84));
	assign Hg72a4 = (~(Efdx84 | Lfdx84));
	assign Tf72a4 = (~(Mv52a4 & Og72a4));
	assign Og72a4 = (Jpnx84 | Huhx84);
	assign Kf62a4 = (Vg72a4 & Ch72a4);
	assign Ch72a4 = (Jh72a4 & Iu42a4);
	assign Jh72a4 = (~(Sc62a4 & Yrbx84));
	assign Sc62a4 = (Nwix84 & Drbx84);
	assign Vg72a4 = (HREADY & Qh72a4);
	assign Qh72a4 = (~(E1dx84 & Ap52a4));
	assign N572a4 = (Me5w84 | HREADY);
	assign Ee4x84 = (!Xh72a4);
	assign Xh72a4 = (HREADY ? Ei72a4 : We62a4);
	assign Ei72a4 = (Li72a4 & Si72a4);
	assign Si72a4 = (~(Zi72a4 & Gj72a4));
	assign Zi72a4 = (Nj72a4 & E7lx84);
	assign Yd4x84 = (!Uj72a4);
	assign Uj72a4 = (HREADY ? Bk72a4 : Mmvx84);
	assign Bk72a4 = (Ik72a4 & Pk72a4);
	assign Pk72a4 = (Wk72a4 & Dl72a4);
	assign Dl72a4 = (Kl72a4 & Rl72a4);
	assign Rl72a4 = (~(W05w84 & Yl72a4));
	assign Yl72a4 = (~(Fm72a4 & Mm72a4));
	assign Mm72a4 = (~(Tm72a4 & An72a4));
	assign An72a4 = (Gf6w84 & Hn72a4);
	assign Hn72a4 = (On72a4 | P0gx84);
	assign Tm72a4 = (Mlbx84 & Gpix84);
	assign Fm72a4 = (Ouhx84 | Xtcx84);
	assign Kl72a4 = (Vn72a4 & Co72a4);
	assign Co72a4 = (~(Jo72a4 & E3ix84));
	assign Jo72a4 = (Gwix84 & Qo72a4);
	assign Qo72a4 = (~(Xo72a4 & Spox84));
	assign Spox84 = (!N052a4);
	assign Xo72a4 = (~(Yrbx84 | N4ix84));
	assign Vn72a4 = (~(Ep72a4 & Atix84));
	assign Ep72a4 = (Lp72a4 & J8cx84);
	assign Lp72a4 = (~(Sp72a4 & Zp72a4));
	assign Zp72a4 = (~(Gq72a4 & Nq72a4));
	assign Nq72a4 = (~(Iokx84 | I86w84));
	assign Gq72a4 = (~(Wcbx84 | Ouhx84));
	assign Sp72a4 = (~(Uq72a4 & X8cx84));
	assign Uq72a4 = (E8dx84 & Br72a4);
	assign Br72a4 = (Nd6w84 | E9cx84);
	assign E9cx84 = (I86w84 & Wcbx84);
	assign Wk72a4 = (Ir72a4 & Pr72a4);
	assign Pr72a4 = (~(Phdx84 & Wr72a4));
	assign Wr72a4 = (~(Ds72a4 & Ks72a4));
	assign Ks72a4 = (~(Xw62a4 & Iqbx84));
	assign Ds72a4 = (Rs72a4 & Ys72a4);
	assign Ys72a4 = (~(Ft72a4 & Hghx84));
	assign Ft72a4 = (Mt72a4 & Wqbx84);
	assign Mt72a4 = (Vvgx84 | Ssex84);
	assign Rs72a4 = (~(Tt72a4 & On72a4));
	assign Tt72a4 = (~(S1dx84 | Pqbx84));
	assign Ir72a4 = (Au72a4 & Hu72a4);
	assign Hu72a4 = (~(Ou72a4 & Pqbx84));
	assign Ou72a4 = (~(J9bx84 & R5cx84));
	assign R5cx84 = (Mzbx84 | Bw2x84);
	assign Au72a4 = (Hgvx84 | T7bx84);
	assign Ik72a4 = (Vu72a4 & Cv72a4);
	assign Cv72a4 = (Jv72a4 & Qv72a4);
	assign Jv72a4 = (Xv72a4 & Ew72a4);
	assign Ew72a4 = (A8ix84 | Yqcx84);
	assign A8ix84 = (!Lowx84);
	assign Lowx84 = (Gwix84 & Lw72a4);
	assign Xv72a4 = (~(Sw72a4 & H6dx84));
	assign Sw72a4 = (~(Zw72a4 & Gx72a4));
	assign Gx72a4 = (Nx72a4 & Ux72a4);
	assign Ux72a4 = (By72a4 & Lncx84);
	assign Lncx84 = (~(Pjwx84 & Huhx84));
	assign Pjwx84 = (C2ix84 & E8dx84);
	assign By72a4 = (Pqix84 & Mtox84);
	assign Mtox84 = (~(Iy72a4 & Ovnx84));
	assign Iy72a4 = (Ggdx84 & Fcdx84);
	assign Ggdx84 = (O8wx84 & Mcdx84);
	assign O8wx84 = (~(R952a4 | Iicx84));
	assign Nx72a4 = (Py72a4 & Wy72a4);
	assign Wy72a4 = (~(Dz72a4 & Yrbx84));
	assign Dz72a4 = (~(W3dx84 | Cuix84));
	assign W3dx84 = (~(Rzhx84 & F2gx84));
	assign Py72a4 = (Kz72a4 & Rz72a4);
	assign Rz72a4 = (~(Yz72a4 & F082a4));
	assign F082a4 = (~(Ba6w84 | Gf6w84));
	assign Yz72a4 = (Xqmx84 & F3mx84);
	assign Xqmx84 = (M082a4 & Evbx84);
	assign M082a4 = (~(N4ix84 | Zg6w84));
	assign Kz72a4 = (~(T082a4 & Zfdx84));
	assign Zfdx84 = (T262a4 & Iicx84);
	assign T082a4 = (Pcbx84 & A182a4);
	assign A182a4 = (~(Ai52a4 & H182a4));
	assign H182a4 = (Ey5w84 | G36w84);
	assign Pcbx84 = (~(Cfcx84 | Iokx84));
	assign Zw72a4 = (O182a4 & V182a4);
	assign V182a4 = (C282a4 & J282a4);
	assign J282a4 = (~(Q282a4 & Qzkx84));
	assign Q282a4 = (~(X282a4 & E382a4));
	assign E382a4 = (~(L382a4 & Ovnx84));
	assign L382a4 = (~(Ifmx84 | Q1xx84));
	assign Ifmx84 = (!Mcdx84);
	assign Mcdx84 = (Tqkx84 & Eobx84);
	assign X282a4 = (~(S382a4 & X8cx84));
	assign X8cx84 = (Ba6w84 & Ub6w84);
	assign S382a4 = (~(Cfcx84 | Efdx84));
	assign C282a4 = (Z382a4 & G482a4);
	assign G482a4 = (~(N482a4 & Soix84));
	assign N482a4 = (~(Ewax84 | N4ix84));
	assign Z382a4 = (~(Fhmx84 & U482a4));
	assign U482a4 = (~(B582a4 & I582a4));
	assign I582a4 = (~(P582a4 & W582a4));
	assign W582a4 = (~(Jfcx84 | Zg6w84));
	assign P582a4 = (Jpnx84 & Ubwx84);
	assign Ubwx84 = (!Efdx84);
	assign B582a4 = (~(D682a4 & X7dx84));
	assign X7dx84 = (K682a4 & Huhx84);
	assign K682a4 = (~(Ba6w84 | Zg6w84));
	assign D682a4 = (Y46w84 & R682a4);
	assign R682a4 = (~(N3cx84 & Y682a4));
	assign Y682a4 = (Z6mx84 | G36w84);
	assign N3cx84 = (Q1xx84 | Ff72a4);
	assign O182a4 = (F782a4 & M782a4);
	assign M782a4 = (Bcix84 | Iokx84);
	assign Bcix84 = (C5mx84 | Ouhx84);
	assign F782a4 = (T782a4 & A882a4);
	assign A882a4 = (~(Mv52a4 & Shix84));
	assign Mv52a4 = (Pcix84 & F3mx84);
	assign T782a4 = (Wd72a4 | Ff72a4);
	assign Ff72a4 = (!N752a4);
	assign N752a4 = (G36w84 & O16w84);
	assign Wd72a4 = (~(H882a4 & Ovnx84));
	assign Ovnx84 = (Oddx84 & Oxlx84);
	assign Oddx84 = (!Cfcx84);
	assign Cfcx84 = (~(O882a4 & F8ox84));
	assign O882a4 = (~(Qtcx84 | Gf6w84));
	assign H882a4 = (~(Efdx84 | Ba6w84));
	assign Efdx84 = (N0mx84 | Wcbx84);
	assign Vu72a4 = (V882a4 & C982a4);
	assign C982a4 = (~(Gc72a4 & J982a4));
	assign V882a4 = (Vx2x84 ? X982a4 : Q982a4);
	assign X982a4 = (Ea82a4 & La82a4);
	assign La82a4 = (~(Gc2y84 & Gwix84));
	assign Gc2y84 = (N4ix84 & Tsix84);
	assign Ea82a4 = (Sa82a4 & Jubx84);
	assign Jubx84 = (!Rfnx84);
	assign Sa82a4 = (~(Za82a4 & Gb82a4));
	assign Gb82a4 = (Nb82a4 & Ub82a4);
	assign Nb82a4 = (~(W05w84 | Hu2x84));
	assign Za82a4 = (Mlbx84 & Plnx84);
	assign Q982a4 = (Mzbx84 | S1dx84);
	assign Sd4x84 = (Wpcx84 ? Bg5w84 : Bc82a4);
	assign Bc82a4 = (~(Qv72a4 & Ic82a4));
	assign Ic82a4 = (~(Pc82a4 & Wc82a4));
	assign Wc82a4 = (~(N4ix84 | D53x84));
	assign Pc82a4 = (~(Dd82a4 | Niix84));
	assign Niix84 = (!Ykwx84);
	assign Dd82a4 = (!Kd82a4);
	assign Qv72a4 = (~(E1dx84 & Lw72a4));
	assign Md4x84 = (~(Rd82a4 & Yd82a4));
	assign Yd82a4 = (Fe82a4 & Mzbx84);
	assign Fe82a4 = (~(J13x84 & Me82a4));
	assign Me82a4 = (~(HREADY & Te82a4));
	assign Te82a4 = (~(Laix84 & Qxmx84));
	assign Rd82a4 = (Af82a4 & Hf82a4);
	assign Hf82a4 = (~(Dt62a4 & A7cx84));
	assign Af82a4 = (~(HREADY & Of82a4));
	assign Of82a4 = (~(Vf82a4 & Cg82a4));
	assign Cg82a4 = (Jg82a4 & Qg82a4);
	assign Qg82a4 = (~(Xg82a4 & W05w84));
	assign Xg82a4 = (Eh82a4 & Qcmx84);
	assign Eh82a4 = (~(Xtcx84 & Lh82a4));
	assign Lh82a4 = (~(Sh82a4 & H6dx84));
	assign Sh82a4 = (~(Zh82a4 & Gi82a4));
	assign Gi82a4 = (~(Hwmx84 & Ewax84));
	assign Zh82a4 = (M6xx84 | Kxcx84);
	assign Jg82a4 = (Ni82a4 & Mg62a4);
	assign Ni82a4 = (~(Ui82a4 & Yybx84));
	assign Ui82a4 = (Tq2x84 & Bj82a4);
	assign Bj82a4 = (~(A0cx84 & Ij82a4));
	assign Ij82a4 = (Fmvx84 | Tsix84);
	assign Vf82a4 = (Pj82a4 & Wj82a4);
	assign Wj82a4 = (~(Nwix84 & Pz2x84));
	assign Pj82a4 = (Dk82a4 & Kk82a4);
	assign Kk82a4 = (~(Rk82a4 & Gwix84));
	assign Rk82a4 = (~(Tsix84 | D53x84));
	assign Dk82a4 = (~(N4ix84 & Yk82a4));
	assign Yk82a4 = (M0px84 | Livx84);
	assign Gd4x84 = (Fl82a4 & Ml82a4);
	assign Ml82a4 = (~(Tl82a4 & Am82a4));
	assign Am82a4 = (Hm82a4 & Om82a4);
	assign Om82a4 = (Vm82a4 & Cn82a4);
	assign Cn82a4 = (Jn82a4 & Pqix84);
	assign Pqix84 = (!Qn82a4);
	assign Jn82a4 = (~(Zymx84 | Y0hx84));
	assign Vm82a4 = (Xn82a4 & Lk52a4);
	assign Lk52a4 = (~(Eo82a4 & Fcdx84));
	assign Eo82a4 = (Uemx84 & Gz4w84);
	assign Xn82a4 = (~(Lo82a4 & Fcdx84));
	assign Lo82a4 = (Benx84 & Ba6w84);
	assign Benx84 = (V1ix84 & Xlkx84);
	assign Hm82a4 = (So82a4 & Zo82a4);
	assign Zo82a4 = (Gp82a4 & Np82a4);
	assign Np82a4 = (~(Up82a4 & L2cx84));
	assign Up82a4 = (Bq82a4 & J8cx84);
	assign Bq82a4 = (~(Iq82a4 & Pq82a4));
	assign Pq82a4 = (Wq82a4 & Dr82a4);
	assign Dr82a4 = (~(Bn42a4 & O16w84));
	assign Wq82a4 = (Kr82a4 & Rr82a4);
	assign Rr82a4 = (~(I86w84 & Yr82a4));
	assign Yr82a4 = (Y46w84 | G9dx84);
	assign Kr82a4 = (Ai52a4 | N0mx84);
	assign N0mx84 = (I86w84 | Y46w84);
	assign Iq82a4 = (S6mx84 & Fs82a4);
	assign Fs82a4 = (Qzkx84 | Wcbx84);
	assign Gp82a4 = (Ms82a4 & Ts82a4);
	assign Ts82a4 = (~(At82a4 & Gwix84));
	assign At82a4 = (Ht82a4 & Hgvx84);
	assign Ht82a4 = (~(Fycx84 & Ot82a4));
	assign Ot82a4 = (~(G4wx84 & E3ix84));
	assign Ms82a4 = (~(Vt82a4 & B9lx84));
	assign Vt82a4 = (~(Tp42a4 | Fn2x84));
	assign So82a4 = (Cu82a4 & Ju82a4);
	assign Ju82a4 = (~(Qu82a4 & Oxlx84));
	assign Qu82a4 = (Gz4w84 & Xu82a4);
	assign Xu82a4 = (~(Ev82a4 & Lv82a4));
	assign Lv82a4 = (~(Ba6w84 & Sv82a4));
	assign Sv82a4 = (~(Zv82a4 & Gw82a4));
	assign Gw82a4 = (Ihdx84 | I86w84);
	assign Zv82a4 = (~(V8wx84 | Ixwx84));
	assign Ev82a4 = (~(Nw82a4 & Xlkx84));
	assign Nw82a4 = (~(Uw82a4 & Bx82a4));
	assign Bx82a4 = (Eobx84 | Iwxx84);
	assign Uw82a4 = (~(Ix82a4 | U3cx84));
	assign Ix82a4 = (Tlwx84 & Px82a4);
	assign Px82a4 = (R952a4 | Iicx84);
	assign Tlwx84 = (I86w84 & Tqkx84);
	assign Cu82a4 = (~(Wx82a4 & W05w84));
	assign Wx82a4 = (Hwmx84 & Ambx84);
	assign Tl82a4 = (Dy82a4 & Ky82a4);
	assign Ky82a4 = (Ry82a4 & Yy82a4);
	assign Yy82a4 = (Fz82a4 & Mz82a4);
	assign Mz82a4 = (~(Gf6w84 & Tz82a4));
	assign Tz82a4 = (~(A092a4 & H092a4));
	assign H092a4 = (Cgix84 | Fcdx84);
	assign Cgix84 = (!Evbx84);
	assign A092a4 = (O092a4 & M172a4);
	assign O092a4 = (E2cx84 | Tqkx84);
	assign Fz82a4 = (V092a4 & C192a4);
	assign C192a4 = (~(Ffox84 & J192a4));
	assign J192a4 = (Pz2x84 | Tq2x84);
	assign V092a4 = (~(Q192a4 & Mmvx84));
	assign Q192a4 = (~(X192a4 & E292a4));
	assign E292a4 = (~(L292a4 & Gc72a4));
	assign L292a4 = (~(Vzcx84 | N4bx84));
	assign X192a4 = (~(S292a4 & Gpbx84));
	assign S292a4 = (~(Z292a4 & G392a4));
	assign G392a4 = (Bdox84 | Fthx84);
	assign Z292a4 = (N392a4 & K5xx84);
	assign K5xx84 = (N4bx84 | Raex84);
	assign Raex84 = (!F2gx84);
	assign N392a4 = (Rybx84 | Tsix84);
	assign Ry82a4 = (U392a4 & B492a4);
	assign B492a4 = (~(V1ix84 & Wn42a4));
	assign Wn42a4 = (Lzlx84 | C2ix84);
	assign U392a4 = (~(Pxbx84 & I492a4));
	assign I492a4 = (~(P492a4 & W492a4));
	assign W492a4 = (D592a4 & K592a4);
	assign K592a4 = (~(R592a4 & Laix84));
	assign R592a4 = (~(Mycx84 | Ulmx84));
	assign D592a4 = (~(Fbex84 | Sbvx84));
	assign P492a4 = (Y592a4 & F692a4);
	assign F692a4 = (~(Hwmx84 & M692a4));
	assign M692a4 = (~(T692a4 & A792a4));
	assign A792a4 = (Ub6w84 | Mw5w84);
	assign Y592a4 = (~(H792a4 & Qxmx84));
	assign H792a4 = (~(Bdox84 & O792a4));
	assign O792a4 = (~(Nacx84 & Vzcx84));
	assign Dy82a4 = (V792a4 & C892a4);
	assign C892a4 = (J892a4 & Q892a4);
	assign Q892a4 = (~(L6mx84 & Uemx84));
	assign J892a4 = (~(Laix84 & A7cx84));
	assign V792a4 = (D072a4 & M6cx84);
	assign M6cx84 = (P1mx84 | H6dx84);
	assign D072a4 = (X892a4 & HREADY);
	assign X892a4 = (E992a4 & Xubx84);
	assign E992a4 = (~(L992a4 & Zo2x84));
	assign L992a4 = (~(V2ox84 | N4ix84));
	assign Fl82a4 = (Fn2x84 | HREADY);
	assign Ad4x84 = (!S992a4);
	assign S992a4 = (Qoox84 ? Z992a4 : Rmnx84);
	assign Z992a4 = (~(Dj0x84 & Vljx84));
	assign Vljx84 = (~(Ga92a4 & Na92a4));
	assign Na92a4 = (Ua92a4 & Bb92a4);
	assign Bb92a4 = (~(Kz0x84 | F11x84));
	assign Ua92a4 = (~(Uv0x84 | Px0x84));
	assign Ga92a4 = (Ib92a4 & Pb92a4);
	assign Pb92a4 = (~(S61x84 | O81x84));
	assign Ib92a4 = (~(A31x84 | W41x84));
	assign Uc4x84 = (!Wb92a4);
	assign Wb92a4 = (HREADY ? Dc92a4 : Wqbx84);
	assign Dc92a4 = (Kc92a4 & Rc92a4);
	assign Rc92a4 = (Yc92a4 & Fd92a4);
	assign Fd92a4 = (Md92a4 & Td92a4);
	assign Td92a4 = (~(Y0hx84 | B9lx84));
	assign Md92a4 = (~(Ejnx84 | Zymx84));
	assign Ejnx84 = (Ae92a4 & Shix84);
	assign Ae92a4 = (~(W05w84 | Nd6w84));
	assign Yc92a4 = (He92a4 & Oe92a4);
	assign Oe92a4 = (~(C2ix84 & Ve92a4));
	assign Ve92a4 = (Evbx84 | Jj52a4);
	assign He92a4 = (Cf92a4 & Jf92a4);
	assign Jf92a4 = (~(Qf92a4 & Wz5w84));
	assign Qf92a4 = (Ey5w84 & Xf92a4);
	assign Xf92a4 = (~(Eg92a4 & Lg92a4));
	assign Lg92a4 = (~(Sg92a4 & Zg92a4));
	assign Zg92a4 = (Gh92a4 & Bn42a4);
	assign Gh92a4 = (S6mx84 & Ub6w84);
	assign Sg92a4 = (Momx84 & Lfdx84);
	assign Lfdx84 = (G36w84 & Jfcx84);
	assign Momx84 = (~(E2cx84 | I86w84));
	assign E2cx84 = (!F8ox84);
	assign Eg92a4 = (~(Nh92a4 & Wcwx84));
	assign Wcwx84 = (C2ix84 & Gz4w84);
	assign Nh92a4 = (~(Ai52a4 | Bhdx84));
	assign Bhdx84 = (!T262a4);
	assign T262a4 = (Uh92a4 & T82y84);
	assign T82y84 = (Bi92a4 & Ii92a4);
	assign Ii92a4 = (Pi92a4 & Sphx84);
	assign Sphx84 = (!Kr5w84);
	assign Pi92a4 = (~(Ct5w84 | Mw5w84));
	assign Bi92a4 = (~(Eobx84 | Tqkx84));
	assign Uh92a4 = (~(Z6mx84 | Uu5w84));
	assign Ai52a4 = (!Ihdx84);
	assign Ihdx84 = (Jfcx84 & Qzkx84);
	assign Cf92a4 = (~(S6mx84 & Wi92a4));
	assign Wi92a4 = (~(C5mx84 & Dj92a4));
	assign Dj92a4 = (~(J5mx84 & Kj92a4));
	assign Kj92a4 = (Rj92a4 | Yj92a4);
	assign Yj92a4 = (Ub6w84 & Fk92a4);
	assign Fk92a4 = (Fcdx84 | Ixwx84);
	assign Rj92a4 = (Y46w84 ? Mk92a4 : Fcdx84);
	assign Mk92a4 = (~(Q1xx84 | Jfcx84));
	assign J5mx84 = (Gz4w84 & J8cx84);
	assign C5mx84 = (~(F8ox84 & J8cx84));
	assign F8ox84 = (Nd6w84 & Gz4w84);
	assign Kc92a4 = (Tk92a4 & Al92a4);
	assign Al92a4 = (Hl92a4 & Ol92a4);
	assign Ol92a4 = (Vl92a4 & Cm92a4);
	assign Cm92a4 = (~(Jm92a4 & Qm92a4));
	assign Qm92a4 = (Xm92a4 | Zvix84);
	assign Vl92a4 = (~(Gwix84 & En92a4));
	assign En92a4 = (Uwix84 | Tn62a4);
	assign Tn62a4 = (~(Vzcx84 | Yqcx84));
	assign Hl92a4 = (Ln92a4 & Sn92a4);
	assign Sn92a4 = (~(Uemx84 & Zn92a4));
	assign Zn92a4 = (~(Go92a4 & No92a4));
	assign No92a4 = (~(Uo92a4 & Tebx84));
	assign Uo92a4 = (~(Bp92a4 & Ip92a4));
	assign Ip92a4 = (~(Pp92a4 & V1ix84));
	assign Pp92a4 = (~(Wcbx84 | Tqkx84));
	assign Bp92a4 = (Zzlx84 | R952a4);
	assign R952a4 = (!Nrnx84);
	assign Go92a4 = (Wp92a4 & F6cx84);
	assign F6cx84 = (!Shix84);
	assign Shix84 = (L2cx84 & Ba6w84);
	assign Wp92a4 = (~(Dq92a4 & G9dx84));
	assign G9dx84 = (!B4cx84);
	assign B4cx84 = (~(Kq92a4 & F1ox84));
	assign Kq92a4 = (~(Qzkx84 | Qklx84));
	assign Qklx84 = (!Uu5w84);
	assign Dq92a4 = (~(Hb52a4 | Zzlx84));
	assign Hb52a4 = (!V8wx84);
	assign Ln92a4 = (~(Pxbx84 & Rq92a4));
	assign Rq92a4 = (~(Yq92a4 & Fr92a4));
	assign Fr92a4 = (Ewax84 | Wqbx84);
	assign Yq92a4 = (Mr92a4 & O8bx84);
	assign Mr92a4 = (~(Gcvx84 & Tr92a4));
	assign Tr92a4 = (Vzcx84 | Xw62a4);
	assign Xw62a4 = (Ulmx84 & Yzhx84);
	assign Ulmx84 = (!Akdx84);
	assign Tk92a4 = (As92a4 & Hs92a4);
	assign Hs92a4 = (Gz4w84 ? Vs92a4 : Os92a4);
	assign Vs92a4 = (Qcmx84 | W05w84);
	assign Os92a4 = (~(Ct92a4 | Jt92a4));
	assign Jt92a4 = (~(Bdox84 | Mmvx84));
	assign Ct92a4 = (Vx2x84 ? U8lx84 : Yevx84);
	assign As92a4 = (Qt92a4 & Xt92a4);
	assign Xt92a4 = (Y4dx84 | Mmvx84);
	assign Qt92a4 = (Xubx84 | Jtcx84);
	assign Xubx84 = (!Symx84);
	assign Symx84 = (W05w84 & Gz4w84);
	assign Oc4x84 = (~(Eu92a4 & Lu92a4));
	assign Lu92a4 = (Su92a4 & Zu92a4);
	assign Zu92a4 = (~(Gv92a4 & Pxbx84));
	assign Gv92a4 = (Sbvx84 & Nv92a4);
	assign Nv92a4 = (Zo2x84 | Kprx84);
	assign Su92a4 = (~(Uv92a4 & S3ix84));
	assign Uv92a4 = (~(Gzfx84 | Gz4w84));
	assign Eu92a4 = (~(Bw92a4 | Iw92a4));
	assign Iw92a4 = (Pw92a4 & J982a4);
	assign Pw92a4 = (~(Ambx84 | Vx2x84));
	assign Bw92a4 = (HREADY ? Ww92a4 : Hu2x84);
	assign Ww92a4 = (~(Dx92a4 & Kx92a4));
	assign Kx92a4 = (Rx92a4 & Yx92a4);
	assign Yx92a4 = (Fy92a4 & My92a4);
	assign My92a4 = (~(Ty92a4 & Az92a4));
	assign Az92a4 = (Lw72a4 | Kd82a4);
	assign Fy92a4 = (Hz92a4 & Oz92a4);
	assign Hz92a4 = (~(Vz92a4 & C0a2a4));
	assign C0a2a4 = (Tp42a4 | W05w84);
	assign Vz92a4 = (J0a2a4 & Qcmx84);
	assign J0a2a4 = (~(Q0a2a4 & Yv42a4));
	assign Q0a2a4 = (~(X0a2a4 & Gpix84));
	assign X0a2a4 = (P0gx84 & Gpbx84);
	assign Rx92a4 = (E1a2a4 & L1a2a4);
	assign L1a2a4 = (~(S1a2a4 & Vvgx84));
	assign Vvgx84 = (!G33x84);
	assign S1a2a4 = (~(Z1a2a4 & G2a2a4));
	assign G2a2a4 = (N2a2a4 & U2a2a4);
	assign U2a2a4 = (Ao62a4 | N4bx84);
	assign N2a2a4 = (B3a2a4 & I3a2a4);
	assign I3a2a4 = (~(P3a2a4 & Ykwx84));
	assign P3a2a4 = (~(Vx2x84 | J13x84));
	assign B3a2a4 = (~(W3a2a4 & B9lx84));
	assign W3a2a4 = (~(Yshx84 | El42a4));
	assign Z1a2a4 = (Dccx84 & D4a2a4);
	assign D4a2a4 = (Yv42a4 | Plnx84);
	assign E1a2a4 = (K4a2a4 & R4a2a4);
	assign R4a2a4 = (~(Rvlx84 & Y4a2a4));
	assign Y4a2a4 = (T0wx84 | F5a2a4);
	assign F5a2a4 = (~(Rybx84 | N4ix84));
	assign K4a2a4 = (~(Pxbx84 & M5a2a4));
	assign M5a2a4 = (~(T5a2a4 & A6a2a4));
	assign A6a2a4 = (~(H6a2a4 & O6a2a4));
	assign O6a2a4 = (~(Ns2x84 | Vx2x84));
	assign H6a2a4 = (~(Akdx84 | Yshx84));
	assign Yshx84 = (!Livx84);
	assign Akdx84 = (Sgcx84 | Tt6w84);
	assign T5a2a4 = (~(V6a2a4 & Fg62a4));
	assign V6a2a4 = (~(Gndx84 & C7a2a4));
	assign C7a2a4 = (Yqcx84 | S1dx84);
	assign Gndx84 = (!Mrcx84);
	assign Dx92a4 = (J7a2a4 & Q7a2a4);
	assign Q7a2a4 = (X7a2a4 & E8a2a4);
	assign X7a2a4 = (L8a2a4 & S8a2a4);
	assign S8a2a4 = (~(Z8a2a4 & H6dx84));
	assign Z8a2a4 = (~(G9a2a4 & N9a2a4));
	assign N9a2a4 = (U9a2a4 & Baa2a4);
	assign Baa2a4 = (~(Iaa2a4 & Bf52a4));
	assign Iaa2a4 = (~(Vzcx84 | Hu2x84));
	assign U9a2a4 = (~(Ty92a4 & Zvix84));
	assign Ty92a4 = (~(Gz4w84 | Pz2x84));
	assign G9a2a4 = (Paa2a4 & Waa2a4);
	assign Waa2a4 = (~(Dba2a4 & J8cx84));
	assign Dba2a4 = (~(M172a4 & Kba2a4));
	assign Kba2a4 = (~(L2cx84 & Rba2a4));
	assign Rba2a4 = (~(Yba2a4 & Fca2a4));
	assign Fca2a4 = (G36w84 | Q66w84);
	assign Yba2a4 = (Mca2a4 & Tca2a4);
	assign Tca2a4 = (~(Ada2a4 & Hda2a4));
	assign Hda2a4 = (~(Oda2a4 & U3cx84));
	assign U3cx84 = (V8wx84 & Wcbx84);
	assign V8wx84 = (I86w84 & Eobx84);
	assign Oda2a4 = (F1ox84 & Uu5w84);
	assign F1ox84 = (Ct5w84 & Kr5w84);
	assign Ada2a4 = (~(Y46w84 & Vda2a4));
	assign Vda2a4 = (Qzkx84 | Tebx84);
	assign Mca2a4 = (Q1xx84 | Jfcx84);
	assign Jfcx84 = (!O16w84);
	assign M172a4 = (!Jj52a4);
	assign Paa2a4 = (Zzlx84 | S6mx84);
	assign S6mx84 = (Gf6w84 & Tqkx84);
	assign Zzlx84 = (!L2cx84);
	assign L8a2a4 = (~(Atix84 & Cea2a4));
	assign Cea2a4 = (~(Jea2a4 & Qea2a4));
	assign Qea2a4 = (Xea2a4 & F3mx84);
	assign Xea2a4 = (~(Efa2a4 & Q1cx84));
	assign Q1cx84 = (!Iwxx84);
	assign Iwxx84 = (Ba6w84 & Wcbx84);
	assign Efa2a4 = (~(Nd6w84 | Gf6w84));
	assign Jea2a4 = (Lfa2a4 & Sfa2a4);
	assign Sfa2a4 = (~(C2ix84 & Zfa2a4));
	assign Zfa2a4 = (~(Gga2a4 & Nga2a4));
	assign Nga2a4 = (Uga2a4 & Z6mx84);
	assign Uga2a4 = (Eobx84 | I86w84);
	assign Gga2a4 = (~(Bha2a4 | Leex84));
	assign Bha2a4 = (G36w84 ? Ixwx84 : Qqmx84);
	assign Qqmx84 = (Q66w84 & Tqkx84);
	assign Lfa2a4 = (Ba6w84 ? Pha2a4 : Iha2a4);
	assign Pha2a4 = (Wha2a4 & Dia2a4);
	assign Dia2a4 = (Nd6w84 ? Ria2a4 : Kia2a4);
	assign Ria2a4 = (C2ix84 | Uemx84);
	assign Kia2a4 = (Q1xx84 | Zg6w84);
	assign Wha2a4 = (Yia2a4 & Fja2a4);
	assign Fja2a4 = (~(Mja2a4 & Xlkx84));
	assign Mja2a4 = (~(Q1xx84 & Z8dx84));
	assign Z8dx84 = (Nrnx84 | I86w84);
	assign Q1xx84 = (!Ixwx84);
	assign Ixwx84 = (Tebx84 & Wcbx84);
	assign Tebx84 = (!I86w84);
	assign Yia2a4 = (Z6mx84 | J8cx84);
	assign Iha2a4 = (~(W8mx84 & Fcdx84));
	assign W8mx84 = (Tja2a4 & Ub6w84);
	assign Tja2a4 = (~(Nd6w84 | Zg6w84));
	assign J7a2a4 = (Aka2a4 & D1gx84);
	assign D1gx84 = (Cubx84 & Hka2a4);
	assign Hka2a4 = (~(Oka2a4 & Vka2a4));
	assign Vka2a4 = (Hwmx84 & Qxmx84);
	assign Oka2a4 = (Mw5w84 & Xgwx84);
	assign Cubx84 = (Mg62a4 | Yybx84);
	assign Aka2a4 = (Vx2x84 ? Jla2a4 : Cla2a4);
	assign Jla2a4 = (Qla2a4 & Xla2a4);
	assign Xla2a4 = (~(E1dx84 & Livx84));
	assign Qla2a4 = (Ema2a4 & Lma2a4);
	assign Lma2a4 = (~(Sma2a4 & Z3px84));
	assign Z3px84 = (~(H8px84 | Gz4w84));
	assign Sma2a4 = (~(Vzcx84 | Kshx84));
	assign Ema2a4 = (~(Y1gx84 & S3ix84));
	assign Cla2a4 = (~(Xgwx84 & Hwmx84));
	assign Xgwx84 = (Plnx84 & Pxbx84);
	assign Ic4x84 = (Gna2a4 ? Zma2a4 : Tc2x84);
	assign Gna2a4 = (Nna2a4 & HREADY);
	assign Zma2a4 = (!HPROT[3]);
	assign Cc4x84 = (Una2a4 ? C92x84 : Nlfx84);
	assign Wb4x84 = (Qoox84 ? Dmux84 : G33x84);
	assign Qb4x84 = (Wpcx84 ? C45w84 : HWRITE);
	assign Kb4x84 = (Wpcx84 ? Ya2x84 : Nna2a4);
	assign Eb4x84 = (~(Boa2a4 & Ioa2a4));
	assign Ioa2a4 = (~(Poa2a4 & HRDATA[31]));
	assign Boa2a4 = (~(G72x84 & Una2a4));
	assign Ya4x84 = (~(Woa2a4 & Dpa2a4));
	assign Dpa2a4 = (~(Poa2a4 & HRDATA[30]));
	assign Woa2a4 = (~(K52x84 & Una2a4));
	assign Sa4x84 = (~(Kpa2a4 & Rpa2a4));
	assign Rpa2a4 = (~(Poa2a4 & HRDATA[29]));
	assign Kpa2a4 = (~(O32x84 & Una2a4));
	assign Ma4x84 = (~(Ypa2a4 & Fqa2a4));
	assign Fqa2a4 = (~(Poa2a4 & HRDATA[28]));
	assign Ypa2a4 = (~(S12x84 & Una2a4));
	assign Ga4x84 = (~(Mqa2a4 & Tqa2a4));
	assign Tqa2a4 = (~(Poa2a4 & HRDATA[27]));
	assign Mqa2a4 = (~(Wz1x84 & Una2a4));
	assign Aa4x84 = (~(Ara2a4 & Hra2a4));
	assign Hra2a4 = (~(Poa2a4 & HRDATA[26]));
	assign Ara2a4 = (~(Ay1x84 & Una2a4));
	assign U94x84 = (~(Ora2a4 & Vra2a4));
	assign Vra2a4 = (~(Poa2a4 & HRDATA[25]));
	assign Ora2a4 = (~(Fw1x84 & Una2a4));
	assign O94x84 = (~(Csa2a4 & Jsa2a4));
	assign Jsa2a4 = (~(Poa2a4 & HRDATA[24]));
	assign Csa2a4 = (~(Ku1x84 & Una2a4));
	assign I94x84 = (~(Qsa2a4 & Xsa2a4));
	assign Xsa2a4 = (~(Poa2a4 & HRDATA[23]));
	assign Qsa2a4 = (~(Ps1x84 & Una2a4));
	assign C94x84 = (~(Eta2a4 & Lta2a4));
	assign Lta2a4 = (~(Poa2a4 & HRDATA[22]));
	assign Eta2a4 = (~(Uq1x84 & Una2a4));
	assign W84x84 = (~(Sta2a4 & Zta2a4));
	assign Zta2a4 = (~(Poa2a4 & HRDATA[21]));
	assign Sta2a4 = (~(Zo1x84 & Una2a4));
	assign Q84x84 = (~(Gua2a4 & Nua2a4));
	assign Nua2a4 = (~(Poa2a4 & HRDATA[20]));
	assign Gua2a4 = (~(En1x84 & Una2a4));
	assign K84x84 = (~(Uua2a4 & Bva2a4));
	assign Bva2a4 = (~(Poa2a4 & HRDATA[19]));
	assign Uua2a4 = (~(Jl1x84 & Una2a4));
	assign E84x84 = (~(Iva2a4 & Pva2a4));
	assign Pva2a4 = (~(Poa2a4 & HRDATA[18]));
	assign Iva2a4 = (~(Oj1x84 & Una2a4));
	assign Y74x84 = (~(Wva2a4 & Dwa2a4));
	assign Dwa2a4 = (~(Poa2a4 & HRDATA[17]));
	assign Wva2a4 = (~(Th1x84 & Una2a4));
	assign S74x84 = (~(Kwa2a4 & Rwa2a4));
	assign Rwa2a4 = (~(Poa2a4 & HRDATA[16]));
	assign Poa2a4 = (~(Nlfx84 | Una2a4));
	assign Kwa2a4 = (~(Yf1x84 & Una2a4));
	assign Una2a4 = (!Crlx84);
	assign M74x84 = (Wpcx84 ? Ig2x84 : Ywa2a4);
	assign Ywa2a4 = (Fxa2a4 & Tplx84);
	assign Fxa2a4 = (Mjkx84 | Bi2x84);
	assign G74x84 = (~(Mxa2a4 & Txa2a4));
	assign Txa2a4 = (~(Aya2a4 & Tplx84));
	assign Aya2a4 = (~(Jrlx84 & Hya2a4));
	assign Hya2a4 = (Wpcx84 | Mjkx84);
	assign Mjkx84 = (!Prax84);
	assign Mxa2a4 = (~(Bi2x84 & Wpcx84));
	assign A74x84 = (H2hx84 ? Oya2a4 : Vs63a4[1]);
	assign U64x84 = (H2hx84 ? Vya2a4 : Vs63a4[0]);
	assign H2hx84 = (HREADY & HPROT[0]);
	assign Vya2a4 = (!Cza2a4);
	assign O64x84 = (~(Jza2a4 & Qza2a4));
	assign Qza2a4 = (~(Xza2a4 & Qdlx84));
	assign Qdlx84 = (E0b2a4 & HREADY);
	assign E0b2a4 = (~(Wnex84 | Pnex84));
	assign Pnex84 = (L0b2a4 & S0b2a4);
	assign S0b2a4 = (Z0b2a4 & Drbx84);
	assign Z0b2a4 = (~(Bw2x84 | J13x84));
	assign L0b2a4 = (G1b2a4 & Aq4w84);
	assign G1b2a4 = (~(B5bx84 | Rybx84));
	assign Wnex84 = (N1b2a4 & U1b2a4);
	assign U1b2a4 = (~(Cavx84 & Ffox84));
	assign N1b2a4 = (Dn52a4 | Ucox84);
	assign Dn52a4 = (~(B2b2a4 & I2b2a4));
	assign B2b2a4 = (~(Rybx84 | Fycx84));
	assign Xza2a4 = (~(W9ex84 | P2b2a4));
	assign P2b2a4 = (Ws4w84 & Lelx84);
	assign Lelx84 = (Cavx84 | Mgnx84);
	assign Jza2a4 = (~(Bh3x84 & Wpcx84));
	assign I64x84 = (~(C64x84 & W2b2a4));
	assign W2b2a4 = (~(D3b2a4 & K3b2a4));
	assign K3b2a4 = (R3b2a4 & Y3b2a4);
	assign Y3b2a4 = (F4b2a4 & M4b2a4);
	assign M4b2a4 = (~(T4b2a4 | HWDATA[30]));
	assign T4b2a4 = (HWDATA[31] | Wz3x84);
	assign F4b2a4 = (~(A5b2a4 | HWDATA[27]));
	assign A5b2a4 = (HWDATA[28] | HWDATA[29]);
	assign R3b2a4 = (H5b2a4 & O5b2a4);
	assign O5b2a4 = (V5b2a4 & HWDATA[26]);
	assign V5b2a4 = (~(Yf1y84 | HWDATA[25]));
	assign H5b2a4 = (~(C6b2a4 | Ezex84));
	assign D3b2a4 = (J6b2a4 & Q6b2a4);
	assign Q6b2a4 = (X6b2a4 & E7b2a4);
	assign E7b2a4 = (L7b2a4 & HWDATA[20]);
	assign L7b2a4 = (~(S7b2a4 | Z7b2a4));
	assign X6b2a4 = (G8b2a4 & N8b2a4);
	assign G8b2a4 = (I6hx84 & Q34x84);
	assign J6b2a4 = (U8b2a4 & B9b2a4);
	assign B9b2a4 = (I9b2a4 & Vhux84);
	assign I9b2a4 = (T14x84 & HWDATA[2]);
	assign U8b2a4 = (Sr0y84 & Lzex84);
	assign Lzex84 = (In4w84 & HWDATA[22]);
	assign Nqax84 = (~(P9b2a4 & W9b2a4));
	assign W9b2a4 = (~(Dab2a4 & D53x84));
	assign Dab2a4 = (Kab2a4 & Ralx84);
	assign Kab2a4 = (~(Rab2a4 & Yab2a4));
	assign Yab2a4 = (~(Fbb2a4 & Mbb2a4));
	assign Mbb2a4 = (~(Tbb2a4 | E7lx84));
	assign Fbb2a4 = (~(Jwgx84 | Hscx84));
	assign Jwgx84 = (!Qoox84);
	assign Qoox84 = (~(Wpcx84 | Ambx84));
	assign Wpcx84 = (!HREADY);
	assign Rab2a4 = (~(Acb2a4 & Nocx84));
	assign Acb2a4 = (~(Ambx84 | V55w84));
	assign P9b2a4 = (~(Uv4w84 & Qwgx84));
	assign Qwgx84 = (~(HREADY & Gz4w84));
	assign Gqax84 = (Ysvx84 ? Axzx84 : Hxzx84);
	assign Zpax84 = (~(Hcb2a4 & Ocb2a4));
	assign Ocb2a4 = (~(Aljx84 & W9ex84));
	assign Hcb2a4 = (Vcb2a4 & Cdb2a4);
	assign Cdb2a4 = (~(HRDATA[4] & S2jx84));
	assign Vcb2a4 = (~(Es0x84 & Enjx84));
	assign Spax84 = (~(Jdb2a4 & Qdb2a4));
	assign Qdb2a4 = (~(Tkjx84 & W9ex84));
	assign Jdb2a4 = (Xdb2a4 & Eeb2a4);
	assign Eeb2a4 = (~(S2jx84 & HRDATA[3]));
	assign Xdb2a4 = (~(Jq0x84 & Enjx84));
	assign Lpax84 = (~(Leb2a4 & Seb2a4));
	assign Seb2a4 = (~(Oo0x84 & Enjx84));
	assign Leb2a4 = (Zeb2a4 & Gfb2a4);
	assign Gfb2a4 = (~(Djjx84 & W9ex84));
	assign Djjx84 = (Nfb2a4 & Ufb2a4);
	assign Nfb2a4 = (Pgb2a4 ? Igb2a4 : Bgb2a4);
	assign Zeb2a4 = (~(S2jx84 & HRDATA[2]));
	assign Epax84 = (~(Wgb2a4 & Dhb2a4));
	assign Dhb2a4 = (~(Pijx84 & W9ex84));
	assign Wgb2a4 = (Khb2a4 & Rhb2a4);
	assign Rhb2a4 = (~(S2jx84 & HRDATA[1]));
	assign Khb2a4 = (~(Tm0x84 & Enjx84));
	assign Xoax84 = (~(Yhb2a4 & Fib2a4));
	assign Fib2a4 = (~(Yjjx84 & W9ex84));
	assign Yhb2a4 = (Mib2a4 & Tib2a4);
	assign Tib2a4 = (~(S2jx84 & HRDATA[0]));
	assign S2jx84 = (Ajb2a4 & F6jx84);
	assign Ajb2a4 = (~(Nlfx84 | X1jx84));
	assign X1jx84 = (!Ulfx84);
	assign Nlfx84 = (~(Hjb2a4 & P25w84));
	assign Hjb2a4 = (~(HRESP | Tc2x84));
	assign Mib2a4 = (~(Yk0x84 & Enjx84));
	assign Enjx84 = (~(Ulfx84 & Ojb2a4));
	assign Ojb2a4 = (W9ex84 | F6jx84);
	assign Ulfx84 = (~(F6jx84 & Vjb2a4));
	assign Vjb2a4 = (~(Ckb2a4 & Jkb2a4));
	assign Jkb2a4 = (~(Jrlx84 | Gz4w84));
	assign Ckb2a4 = (Crlx84 & Prax84);
	assign Crlx84 = (Ya2x84 & HREADY);
	assign F6jx84 = (~(W9ex84 | Dj0x84));
	assign W9ex84 = (~(Li72a4 & Qkb2a4));
	assign Qkb2a4 = (~(Xkb2a4 & Elb2a4));
	assign Elb2a4 = (~(Llb2a4 | Kehx84));
	assign Kehx84 = (Ffhx84 & Nr4w84);
	assign Ffhx84 = (Slb2a4 & Zlb2a4);
	assign Zlb2a4 = (~(Gmb2a4 & Ap6w84));
	assign Gmb2a4 = (P7gx84 & Bf0y84);
	assign Llb2a4 = (~(Nj72a4 & E7lx84));
	assign Xkb2a4 = (Nmb2a4 & Umb2a4);
	assign Umb2a4 = (Slb2a4 | Oghx84);
	assign Slb2a4 = (~(Bnb2a4 & Inb2a4));
	assign Inb2a4 = (Pnb2a4 & Wnb2a4);
	assign Wnb2a4 = (~(Dob2a4 & F1vx84));
	assign F1vx84 = (Kob2a4 & Rob2a4);
	assign Rob2a4 = (Kkbx84 | Pzux84);
	assign Pzux84 = (Yob2a4 & Fpb2a4);
	assign Fpb2a4 = (Mpb2a4 & Tpb2a4);
	assign Tpb2a4 = (~(Aqb2a4 & Nr62a4));
	assign Aqb2a4 = (~(Pqbx84 | Zo2x84));
	assign Mpb2a4 = (~(Wyox84 | Vwfx84));
	assign Vwfx84 = (~(Ivrx84 | Gz4w84));
	assign Ivrx84 = (Sbox84 | B5bx84);
	assign Yob2a4 = (Hqb2a4 & Oqb2a4);
	assign Oqb2a4 = (~(Gz4w84 & Vqb2a4));
	assign Vqb2a4 = (~(Crb2a4 & Jrb2a4));
	assign Jrb2a4 = (Qrb2a4 & Xrb2a4);
	assign Xrb2a4 = (Cuix84 | Fn2x84);
	assign Qrb2a4 = (Uy1y84 | Bw2x84);
	assign Crb2a4 = (Esb2a4 & Lsb2a4);
	assign Lsb2a4 = (Tswx84 | Tq2x84);
	assign Esb2a4 = (B5bx84 | Evix84);
	assign Hqb2a4 = (Hu2x84 ? Zsb2a4 : Ssb2a4);
	assign Zsb2a4 = (~(Zvix84 & Ambx84));
	assign Ssb2a4 = (Bs1y84 | Wbcx84);
	assign Kob2a4 = (Oghx84 | Gyux84);
	assign Gyux84 = (Gtb2a4 & Ntb2a4);
	assign Ntb2a4 = (~(L3ix84 & A2ox84));
	assign Gtb2a4 = (Utb2a4 & Bub2a4);
	assign Bub2a4 = (~(Iub2a4 & Devx84));
	assign Devx84 = (~(Fn2x84 | Vx2x84));
	assign Iub2a4 = (~(Xtcx84 | Evix84));
	assign Utb2a4 = (~(Pub2a4 & H6dx84));
	assign Pub2a4 = (~(Wub2a4 & Dvb2a4));
	assign Dvb2a4 = (~(Kvb2a4 & U8lx84));
	assign Kvb2a4 = (~(Ucox84 | Wqbx84));
	assign Wub2a4 = (~(Rvb2a4 & Gpix84));
	assign Rvb2a4 = (~(Evix84 | Pz2x84));
	assign Dob2a4 = (M1vx84 & Y0vx84);
	assign Y0vx84 = (Yvb2a4 | Izux84);
	assign Izux84 = (Fwb2a4 & Mwb2a4);
	assign Mwb2a4 = (Twb2a4 & L42y84);
	assign L42y84 = (Axb2a4 & Hxb2a4);
	assign Hxb2a4 = (~(Oxb2a4 & Gpix84));
	assign Oxb2a4 = (~(Fmvx84 | Hgvx84));
	assign Twb2a4 = (Vxb2a4 & Cyb2a4);
	assign Cyb2a4 = (~(Jyb2a4 & Yqcx84));
	assign Jyb2a4 = (~(Bw2x84 | Pz2x84));
	assign Vxb2a4 = (~(Yevx84 & Yzhx84));
	assign Yevx84 = (Hu2x84 & Mmvx84);
	assign Fwb2a4 = (~(Qyb2a4 | Xyb2a4));
	assign Xyb2a4 = (J13x84 ? F352a4 : Ezb2a4);
	assign Ezb2a4 = (~(Lzb2a4 & Szb2a4));
	assign Szb2a4 = (Vx2x84 | Pz2x84);
	assign Lzb2a4 = (~(Zzb2a4 | Jq52a4));
	assign Zzb2a4 = (~(Quix84 | Mmvx84));
	assign Quix84 = (!G0c2a4);
	assign Qyb2a4 = (~(N0c2a4 & U0c2a4));
	assign U0c2a4 = (Hu2x84 ? B1c2a4 : Naxx84);
	assign N0c2a4 = (Ns2x84 ? P1c2a4 : I1c2a4);
	assign P1c2a4 = (W1c2a4 | Wbcx84);
	assign I1c2a4 = (D2c2a4 & Xw1y84);
	assign Xw1y84 = (Rybx84 | Hu2x84);
	assign D2c2a4 = (K2c2a4 & Ambx84);
	assign M1vx84 = (R2c2a4 & Y2c2a4);
	assign Y2c2a4 = (B0gx84 | Bw2x84);
	assign R2c2a4 = (~(Tu1y84 | Ws62a4));
	assign Ws62a4 = (Pxbx84 & Pqbx84);
	assign Tu1y84 = (F3c2a4 & J13x84);
	assign F3c2a4 = (~(A2ox84 | F352a4));
	assign Pnb2a4 = (~(N4ix84 | Ns2x84));
	assign Bnb2a4 = (~(W1c2a4 | Wbcx84));
	assign Nmb2a4 = (Gj72a4 & M3c2a4);
	assign M3c2a4 = (~(T3c2a4 & A4c2a4));
	assign A4c2a4 = (~(Yn0y84 | Wl6w84));
	assign T3c2a4 = (Ap6w84 & P7gx84);
	assign P7gx84 = (~(H4c2a4 & O4c2a4));
	assign O4c2a4 = (~(V4c2a4 & Qxmx84));
	assign H4c2a4 = (Mzbx84 | P1mx84);
	assign Gj72a4 = (~(C5c2a4 & J5c2a4));
	assign J5c2a4 = (Q5c2a4 | X5c2a4);
	assign X5c2a4 = (Pgb2a4 ? L6c2a4 : E6c2a4);
	assign Q5c2a4 = (~(S6c2a4 & Z6c2a4));
	assign S6c2a4 = (~(G7c2a4 & N7c2a4));
	assign N7c2a4 = (U7c2a4 | B8c2a4);
	assign C5c2a4 = (I8c2a4 & P8c2a4);
	assign I8c2a4 = (W8c2a4 | B8c2a4);
	assign B8c2a4 = (Pgb2a4 & D9c2a4);
	assign W8c2a4 = (U7c2a4 | G7c2a4);
	assign U7c2a4 = (K9c2a4 & R9c2a4);
	assign Li72a4 = (~(Y9c2a4 & Cwgx84));
	assign Cwgx84 = (!Ilux84);
	assign Ilux84 = (Dmux84 & Tbb2a4);
	assign Y9c2a4 = (~(Mhfx84 & Fac2a4));
	assign Fac2a4 = (Mac2a4 | Dmux84);
	assign Mac2a4 = (!Cc3x84);
	assign Qoax84 = (~(Tac2a4 & Abc2a4));
	assign Abc2a4 = (~(Cx8w84 & L0ex84));
	assign Tac2a4 = (Hbc2a4 & Obc2a4);
	assign Obc2a4 = (~(Jzdx84 & Vbc2a4));
	assign Vbc2a4 = (~(Cza2a4 & Ccc2a4));
	assign Ccc2a4 = (~(P25w84 & Jcc2a4));
	assign Jcc2a4 = (~(Jnwx84 & Qcc2a4));
	assign Qcc2a4 = (~(Jpnx84 & Bn42a4));
	assign Jpnx84 = (V1ix84 & Tqkx84);
	assign V1ix84 = (~(Gpbx84 | Nd6w84));
	assign Jnwx84 = (!L6mx84);
	assign Hbc2a4 = (~(Czdx84 & Nj63a4[0]));
	assign Czdx84 = (Xcc2a4 & Edc2a4);
	assign Xcc2a4 = (~(Ambx84 | Pz2x84));
	assign Joax84 = (~(Ldc2a4 & Sdc2a4));
	assign Sdc2a4 = (~(Y79w84 & L0ex84));
	assign Ldc2a4 = (Zdc2a4 & Gec2a4);
	assign Gec2a4 = (~(Jzdx84 & HADDR[6]));
	assign Zdc2a4 = (~(Tk63a4[5] & E0ex84));
	assign Coax84 = (~(Nec2a4 & Uec2a4));
	assign Uec2a4 = (~(T99w84 & L0ex84));
	assign Nec2a4 = (Bfc2a4 & Ifc2a4);
	assign Ifc2a4 = (~(Jzdx84 & HADDR[7]));
	assign Bfc2a4 = (~(Tk63a4[6] & E0ex84));
	assign Vnax84 = (~(Pfc2a4 & Wfc2a4));
	assign Wfc2a4 = (~(Ob9w84 & L0ex84));
	assign Pfc2a4 = (Dgc2a4 & Kgc2a4);
	assign Kgc2a4 = (~(Jzdx84 & HADDR[8]));
	assign Dgc2a4 = (~(Tk63a4[7] & E0ex84));
	assign Onax84 = (~(Rgc2a4 & Ygc2a4));
	assign Ygc2a4 = (~(Ef9w84 & L0ex84));
	assign Rgc2a4 = (Fhc2a4 & Mhc2a4);
	assign Mhc2a4 = (~(Jzdx84 & HADDR[10]));
	assign Fhc2a4 = (~(Tk63a4[9] & E0ex84));
	assign Hnax84 = (~(Thc2a4 & Aic2a4));
	assign Aic2a4 = (~(Ah9w84 & L0ex84));
	assign Thc2a4 = (Hic2a4 & Oic2a4);
	assign Oic2a4 = (~(Jzdx84 & HADDR[11]));
	assign Hic2a4 = (~(Tk63a4[10] & E0ex84));
	assign Anax84 = (~(Vic2a4 & Cjc2a4));
	assign Cjc2a4 = (~(Wi9w84 & L0ex84));
	assign Vic2a4 = (Jjc2a4 & Qjc2a4);
	assign Qjc2a4 = (~(Jzdx84 & HADDR[12]));
	assign Jjc2a4 = (~(Tk63a4[11] & E0ex84));
	assign Tmax84 = (~(Xjc2a4 & Ekc2a4));
	assign Ekc2a4 = (~(Sk9w84 & L0ex84));
	assign Xjc2a4 = (Lkc2a4 & Skc2a4);
	assign Skc2a4 = (~(Jzdx84 & HADDR[13]));
	assign Lkc2a4 = (~(Tk63a4[12] & E0ex84));
	assign Mmax84 = (~(Zkc2a4 & Glc2a4));
	assign Glc2a4 = (~(Om9w84 & L0ex84));
	assign Zkc2a4 = (Nlc2a4 & Ulc2a4);
	assign Ulc2a4 = (~(Jzdx84 & HADDR[14]));
	assign Nlc2a4 = (~(Tk63a4[13] & E0ex84));
	assign Fmax84 = (~(Bmc2a4 & Imc2a4));
	assign Imc2a4 = (~(Ko9w84 & L0ex84));
	assign Bmc2a4 = (Pmc2a4 & Wmc2a4);
	assign Wmc2a4 = (~(Jzdx84 & HADDR[15]));
	assign Pmc2a4 = (~(Tk63a4[14] & E0ex84));
	assign Ylax84 = (~(Dnc2a4 & Knc2a4));
	assign Knc2a4 = (~(Gq9w84 & L0ex84));
	assign Dnc2a4 = (Rnc2a4 & Ync2a4);
	assign Ync2a4 = (~(Jzdx84 & HADDR[16]));
	assign Rnc2a4 = (~(Tk63a4[15] & E0ex84));
	assign Rlax84 = (~(Foc2a4 & Moc2a4));
	assign Moc2a4 = (~(Cs9w84 & L0ex84));
	assign Foc2a4 = (Toc2a4 & Apc2a4);
	assign Apc2a4 = (~(Jzdx84 & HADDR[17]));
	assign Toc2a4 = (~(Tk63a4[16] & E0ex84));
	assign Klax84 = (~(Hpc2a4 & Opc2a4));
	assign Opc2a4 = (~(Yt9w84 & L0ex84));
	assign Hpc2a4 = (Vpc2a4 & Cqc2a4);
	assign Cqc2a4 = (~(Jzdx84 & HADDR[18]));
	assign Vpc2a4 = (~(Tk63a4[17] & E0ex84));
	assign Dlax84 = (~(Jqc2a4 & Qqc2a4));
	assign Qqc2a4 = (~(Uv9w84 & L0ex84));
	assign Jqc2a4 = (Xqc2a4 & Erc2a4);
	assign Erc2a4 = (~(Jzdx84 & HADDR[19]));
	assign Xqc2a4 = (~(Tk63a4[18] & E0ex84));
	assign Wkax84 = (~(Lrc2a4 & Src2a4));
	assign Src2a4 = (~(Qx9w84 & L0ex84));
	assign Lrc2a4 = (Zrc2a4 & Gsc2a4);
	assign Gsc2a4 = (~(Jzdx84 & HADDR[20]));
	assign Zrc2a4 = (~(Tk63a4[19] & E0ex84));
	assign Pkax84 = (~(Nsc2a4 & Usc2a4));
	assign Usc2a4 = (~(Mz9w84 & L0ex84));
	assign Nsc2a4 = (Btc2a4 & Itc2a4);
	assign Itc2a4 = (~(Jzdx84 & HADDR[21]));
	assign Btc2a4 = (~(Tk63a4[20] & E0ex84));
	assign Ikax84 = (~(Ptc2a4 & Wtc2a4));
	assign Wtc2a4 = (~(I1aw84 & L0ex84));
	assign Ptc2a4 = (Duc2a4 & Kuc2a4);
	assign Kuc2a4 = (~(Jzdx84 & HADDR[22]));
	assign Duc2a4 = (~(Tk63a4[21] & E0ex84));
	assign Bkax84 = (~(Ruc2a4 & Yuc2a4));
	assign Yuc2a4 = (~(E3aw84 & L0ex84));
	assign Ruc2a4 = (Fvc2a4 & Mvc2a4);
	assign Mvc2a4 = (~(Jzdx84 & HADDR[23]));
	assign Fvc2a4 = (~(Tk63a4[22] & E0ex84));
	assign Ujax84 = (~(Tvc2a4 & Awc2a4));
	assign Awc2a4 = (~(W6aw84 & L0ex84));
	assign Tvc2a4 = (Hwc2a4 & Owc2a4);
	assign Owc2a4 = (~(Jzdx84 & HADDR[25]));
	assign Hwc2a4 = (~(Tk63a4[24] & E0ex84));
	assign Njax84 = (~(Vwc2a4 & Cxc2a4));
	assign Cxc2a4 = (~(S8aw84 & L0ex84));
	assign Vwc2a4 = (Jxc2a4 & Qxc2a4);
	assign Qxc2a4 = (~(Jzdx84 & HADDR[26]));
	assign Jxc2a4 = (~(Tk63a4[25] & E0ex84));
	assign Gjax84 = (~(Xxc2a4 & Eyc2a4));
	assign Eyc2a4 = (~(Oaaw84 & L0ex84));
	assign Xxc2a4 = (Lyc2a4 & Syc2a4);
	assign Syc2a4 = (~(Jzdx84 & HADDR[27]));
	assign Jzdx84 = (Edc2a4 & Zyc2a4);
	assign Zyc2a4 = (~(Gzc2a4 & Nzc2a4));
	assign Nzc2a4 = (Jxmx84 | Pqbx84);
	assign Gzc2a4 = (Uzc2a4 & Fmvx84);
	assign Uzc2a4 = (~(B0d2a4 & Ambx84));
	assign B0d2a4 = (~(Gwbx84 & J8cx84));
	assign Edc2a4 = (!L0ex84);
	assign Lyc2a4 = (~(Tk63a4[26] & E0ex84));
	assign E0ex84 = (~(L0ex84 | J9bx84));
	assign L0ex84 = (~(HREADY & I0d2a4));
	assign I0d2a4 = (~(P0d2a4 & W0d2a4));
	assign W0d2a4 = (D1d2a4 & K1d2a4);
	assign K1d2a4 = (R1d2a4 & Y1d2a4);
	assign R1d2a4 = (Oz92a4 & Qnix84);
	assign Oz92a4 = (~(F2d2a4 & Hbmx84));
	assign Hbmx84 = (Qvax84 & Tsix84);
	assign F2d2a4 = (~(Zo2x84 | Hu2x84));
	assign D1d2a4 = (M2d2a4 & T2d2a4);
	assign T2d2a4 = (~(A3d2a4 & Jj52a4));
	assign Jj52a4 = (L2cx84 & Nd6w84);
	assign A3d2a4 = (~(L4ox84 | Qtcx84));
	assign L4ox84 = (!Lzlx84);
	assign Lzlx84 = (Zg6w84 & Tqkx84);
	assign Tqkx84 = (!Ba6w84);
	assign M2d2a4 = (H3d2a4 & O3d2a4);
	assign O3d2a4 = (~(V3d2a4 & C4d2a4));
	assign C4d2a4 = (~(Gpbx84 | Ba6w84));
	assign V3d2a4 = (Fhmx84 & Oxlx84);
	assign H3d2a4 = (~(J4d2a4 & Rzhx84));
	assign J4d2a4 = (~(Naxx84 | H8px84));
	assign Naxx84 = (!Ghxx84);
	assign Ghxx84 = (Yzhx84 & Yqcx84);
	assign P0d2a4 = (Q4d2a4 & X4d2a4);
	assign X4d2a4 = (E5d2a4 & L5d2a4);
	assign L5d2a4 = (~(Wadx84 & Z6mx84));
	assign Z6mx84 = (!Fcdx84);
	assign Fcdx84 = (I86w84 & Q66w84);
	assign Wadx84 = (Evbx84 & Edmx84);
	assign Evbx84 = (L6mx84 & Leex84);
	assign L6mx84 = (Ub6w84 & Gz4w84);
	assign E5d2a4 = (S5d2a4 & Z5d2a4);
	assign Z5d2a4 = (Wjwx84 | G6d2a4);
	assign G6d2a4 = (Gwbx84 & N6d2a4);
	assign N6d2a4 = (~(Bn42a4 & Nrnx84));
	assign Bn42a4 = (~(Eobx84 | Wcbx84));
	assign Wcbx84 = (!Q66w84);
	assign Eobx84 = (!Y46w84);
	assign Gwbx84 = (~(I86w84 | Ba6w84));
	assign Wjwx84 = (~(U6d2a4 & Uemx84));
	assign Uemx84 = (Gf6w84 & J8cx84);
	assign U6d2a4 = (Huhx84 & E8dx84);
	assign Huhx84 = (L2cx84 & Leex84);
	assign Leex84 = (!Nd6w84);
	assign L2cx84 = (Gz4w84 & Iokx84);
	assign S5d2a4 = (~(Phdx84 & B7d2a4));
	assign B7d2a4 = (Dzox84 | Jq52a4);
	assign Jq52a4 = (Hghx84 & Gcvx84);
	assign Q4d2a4 = (I7d2a4 & P7d2a4);
	assign I7d2a4 = (W7d2a4 & D8d2a4);
	assign D8d2a4 = (~(Frcx84 & Rfnx84));
	assign Rfnx84 = (Gwix84 & Tq2x84);
	assign W7d2a4 = (Gqox84 | Jxmx84);
	assign Ziax84 = (~(K8d2a4 & R8d2a4));
	assign R8d2a4 = (~(Y8d2a4 & Pu63a4[23]));
	assign K8d2a4 = (F9d2a4 & M9d2a4);
	assign M9d2a4 = (~(T9d2a4 & X473a4[23]));
	assign F9d2a4 = (~(H173a4[23] & Aad2a4));
	assign Siax84 = (~(Had2a4 & Oad2a4));
	assign Oad2a4 = (~(Y8d2a4 & Pu63a4[22]));
	assign Had2a4 = (Vad2a4 & Cbd2a4);
	assign Cbd2a4 = (~(T9d2a4 & X473a4[22]));
	assign Vad2a4 = (~(H173a4[22] & Aad2a4));
	assign Liax84 = (~(Jbd2a4 & Qbd2a4));
	assign Qbd2a4 = (~(Y8d2a4 & Pu63a4[21]));
	assign Jbd2a4 = (Xbd2a4 & Ecd2a4);
	assign Ecd2a4 = (~(T9d2a4 & X473a4[21]));
	assign Xbd2a4 = (~(H173a4[21] & Aad2a4));
	assign Eiax84 = (~(Lcd2a4 & Scd2a4));
	assign Scd2a4 = (~(Y8d2a4 & Pu63a4[20]));
	assign Lcd2a4 = (Zcd2a4 & Gdd2a4);
	assign Gdd2a4 = (~(T9d2a4 & X473a4[20]));
	assign Zcd2a4 = (~(H173a4[20] & Aad2a4));
	assign Xhax84 = (~(Ndd2a4 & Udd2a4));
	assign Udd2a4 = (~(Y8d2a4 & Pu63a4[19]));
	assign Ndd2a4 = (Bed2a4 & Ied2a4);
	assign Ied2a4 = (~(T9d2a4 & X473a4[19]));
	assign Bed2a4 = (~(H173a4[19] & Aad2a4));
	assign Qhax84 = (~(Ped2a4 & Wed2a4));
	assign Wed2a4 = (~(Y8d2a4 & Pu63a4[18]));
	assign Ped2a4 = (Dfd2a4 & Kfd2a4);
	assign Kfd2a4 = (~(T9d2a4 & X473a4[18]));
	assign Dfd2a4 = (~(H173a4[18] & Aad2a4));
	assign Jhax84 = (~(Rfd2a4 & Yfd2a4));
	assign Yfd2a4 = (~(Y8d2a4 & Pu63a4[17]));
	assign Rfd2a4 = (Fgd2a4 & Mgd2a4);
	assign Mgd2a4 = (~(T9d2a4 & X473a4[17]));
	assign Fgd2a4 = (~(H173a4[17] & Aad2a4));
	assign Chax84 = (~(Tgd2a4 & Ahd2a4));
	assign Ahd2a4 = (~(Y8d2a4 & Pu63a4[16]));
	assign Tgd2a4 = (Hhd2a4 & Ohd2a4);
	assign Ohd2a4 = (~(T9d2a4 & X473a4[16]));
	assign Hhd2a4 = (~(H173a4[16] & Aad2a4));
	assign Vgax84 = (~(Vhd2a4 & Cid2a4));
	assign Cid2a4 = (~(Y8d2a4 & Pu63a4[15]));
	assign Vhd2a4 = (Jid2a4 & Qid2a4);
	assign Qid2a4 = (~(T9d2a4 & X473a4[15]));
	assign Jid2a4 = (~(H173a4[15] & Aad2a4));
	assign Ogax84 = (~(Xid2a4 & Ejd2a4));
	assign Ejd2a4 = (~(Y8d2a4 & Pu63a4[14]));
	assign Xid2a4 = (Ljd2a4 & Sjd2a4);
	assign Sjd2a4 = (~(T9d2a4 & X473a4[14]));
	assign Ljd2a4 = (~(H173a4[14] & Aad2a4));
	assign Hgax84 = (~(Zjd2a4 & Gkd2a4));
	assign Gkd2a4 = (~(Y8d2a4 & Pu63a4[13]));
	assign Zjd2a4 = (Nkd2a4 & Ukd2a4);
	assign Ukd2a4 = (~(T9d2a4 & X473a4[13]));
	assign Nkd2a4 = (~(H173a4[13] & Aad2a4));
	assign Agax84 = (~(Bld2a4 & Ild2a4));
	assign Ild2a4 = (~(Y8d2a4 & Pu63a4[12]));
	assign Bld2a4 = (Pld2a4 & Wld2a4);
	assign Wld2a4 = (~(T9d2a4 & X473a4[12]));
	assign Pld2a4 = (~(H173a4[12] & Aad2a4));
	assign Tfax84 = (~(Dmd2a4 & Kmd2a4));
	assign Kmd2a4 = (~(Y8d2a4 & Pu63a4[11]));
	assign Dmd2a4 = (Rmd2a4 & Ymd2a4);
	assign Ymd2a4 = (~(T9d2a4 & X473a4[11]));
	assign Rmd2a4 = (~(H173a4[11] & Aad2a4));
	assign Mfax84 = (~(Fnd2a4 & Mnd2a4));
	assign Mnd2a4 = (~(Y8d2a4 & Pu63a4[10]));
	assign Fnd2a4 = (Tnd2a4 & Aod2a4);
	assign Aod2a4 = (~(T9d2a4 & X473a4[10]));
	assign Tnd2a4 = (~(H173a4[10] & Aad2a4));
	assign Ffax84 = (~(Hod2a4 & Ood2a4));
	assign Ood2a4 = (~(Y8d2a4 & Pu63a4[9]));
	assign Hod2a4 = (Vod2a4 & Cpd2a4);
	assign Cpd2a4 = (~(T9d2a4 & X473a4[9]));
	assign Vod2a4 = (~(H173a4[9] & Aad2a4));
	assign Yeax84 = (~(Jpd2a4 & Qpd2a4));
	assign Qpd2a4 = (~(Y8d2a4 & Pu63a4[8]));
	assign Jpd2a4 = (Xpd2a4 & Eqd2a4);
	assign Eqd2a4 = (~(T9d2a4 & X473a4[8]));
	assign Xpd2a4 = (~(H173a4[8] & Aad2a4));
	assign Reax84 = (~(Lqd2a4 & Sqd2a4));
	assign Sqd2a4 = (~(Y8d2a4 & Pu63a4[7]));
	assign Lqd2a4 = (Zqd2a4 & Grd2a4);
	assign Grd2a4 = (~(T9d2a4 & X473a4[7]));
	assign Zqd2a4 = (~(H173a4[7] & Aad2a4));
	assign Keax84 = (~(Nrd2a4 & Urd2a4));
	assign Urd2a4 = (~(Y8d2a4 & Pu63a4[6]));
	assign Nrd2a4 = (Bsd2a4 & Isd2a4);
	assign Isd2a4 = (~(T9d2a4 & X473a4[6]));
	assign Bsd2a4 = (~(H173a4[6] & Aad2a4));
	assign Deax84 = (~(Psd2a4 & Wsd2a4));
	assign Wsd2a4 = (~(Y8d2a4 & Pu63a4[5]));
	assign Psd2a4 = (Dtd2a4 & Ktd2a4);
	assign Ktd2a4 = (~(T9d2a4 & X473a4[5]));
	assign Dtd2a4 = (~(H173a4[5] & Aad2a4));
	assign Wdax84 = (~(Rtd2a4 & Ytd2a4));
	assign Ytd2a4 = (~(Y8d2a4 & Pu63a4[4]));
	assign Rtd2a4 = (Fud2a4 & Mud2a4);
	assign Mud2a4 = (~(T9d2a4 & X473a4[4]));
	assign Fud2a4 = (~(H173a4[4] & Aad2a4));
	assign Pdax84 = (~(Tud2a4 & Avd2a4));
	assign Avd2a4 = (~(Y8d2a4 & Pu63a4[3]));
	assign Tud2a4 = (Hvd2a4 & Ovd2a4);
	assign Ovd2a4 = (~(T9d2a4 & X473a4[3]));
	assign Hvd2a4 = (~(H173a4[3] & Aad2a4));
	assign Idax84 = (~(Vvd2a4 & Cwd2a4));
	assign Cwd2a4 = (~(Y8d2a4 & Pu63a4[2]));
	assign Vvd2a4 = (Jwd2a4 & Qwd2a4);
	assign Qwd2a4 = (~(T9d2a4 & X473a4[2]));
	assign Jwd2a4 = (~(H173a4[2] & Aad2a4));
	assign Bdax84 = (~(Xwd2a4 & Exd2a4));
	assign Exd2a4 = (~(Y8d2a4 & Pu63a4[1]));
	assign Xwd2a4 = (Lxd2a4 & Sxd2a4);
	assign Sxd2a4 = (~(T9d2a4 & X473a4[1]));
	assign Lxd2a4 = (~(H173a4[1] & Aad2a4));
	assign Ucax84 = (~(Zxd2a4 & Gyd2a4));
	assign Gyd2a4 = (~(Y8d2a4 & Pu63a4[0]));
	assign Zxd2a4 = (Nyd2a4 & Uyd2a4);
	assign Uyd2a4 = (~(T9d2a4 & X473a4[0]));
	assign T9d2a4 = (Bzd2a4 & Izd2a4);
	assign Bzd2a4 = (~(Y8d2a4 | Nchx84));
	assign Nyd2a4 = (~(H173a4[0] & Aad2a4));
	assign Aad2a4 = (~(Pzd2a4 | Izd2a4));
	assign Izd2a4 = (Pdhx84 & Wzd2a4);
	assign Wzd2a4 = (!Pu63a4[0]);
	assign Pdhx84 = (D0e2a4 & K0e2a4);
	assign K0e2a4 = (R0e2a4 & Y0e2a4);
	assign Y0e2a4 = (F1e2a4 & M1e2a4);
	assign M1e2a4 = (~(T1e2a4 | Pu63a4[7]));
	assign T1e2a4 = (Pu63a4[8] | Pu63a4[9]);
	assign F1e2a4 = (~(A2e2a4 | Pu63a4[4]));
	assign A2e2a4 = (Pu63a4[5] | Pu63a4[6]);
	assign R0e2a4 = (H2e2a4 & O2e2a4);
	assign O2e2a4 = (~(V2e2a4 | Pu63a4[23]));
	assign V2e2a4 = (Pu63a4[2] | Pu63a4[3]);
	assign H2e2a4 = (~(C3e2a4 | Pu63a4[20]));
	assign C3e2a4 = (Pu63a4[21] | Pu63a4[22]);
	assign D0e2a4 = (J3e2a4 & Q3e2a4);
	assign Q3e2a4 = (X3e2a4 & E4e2a4);
	assign E4e2a4 = (~(L4e2a4 | Pu63a4[18]));
	assign L4e2a4 = (Pu63a4[19] | Pu63a4[1]);
	assign X3e2a4 = (~(S4e2a4 | Pu63a4[15]));
	assign S4e2a4 = (Pu63a4[16] | Pu63a4[17]);
	assign J3e2a4 = (Z4e2a4 & G5e2a4);
	assign G5e2a4 = (~(N5e2a4 | Pu63a4[12]));
	assign N5e2a4 = (Pu63a4[13] | Pu63a4[14]);
	assign Z4e2a4 = (~(Pu63a4[10] | Pu63a4[11]));
	assign Pzd2a4 = (Y8d2a4 | Nchx84);
	assign Y8d2a4 = (~(Idhx84 | Nchx84));
	assign Nchx84 = (U5e2a4 & B6e2a4);
	assign B6e2a4 = (Ebhx84 & In4w84);
	assign Ebhx84 = (~(Dfgx84 | Q34x84));
	assign U5e2a4 = (R7hx84 & T14x84);
	assign Idhx84 = (Mq3x84 & I6e2a4);
	assign I6e2a4 = (STCLKEN | P6e2a4);
	assign Ncax84 = (~(W6e2a4 & D7e2a4));
	assign D7e2a4 = (K7e2a4 | Nocx84);
	assign W6e2a4 = (R7e2a4 & Y7e2a4);
	assign Y7e2a4 = (F8e2a4 | Tmhx84);
	assign Tmhx84 = (M8e2a4 & T8e2a4);
	assign T8e2a4 = (A9e2a4 & H9e2a4);
	assign H9e2a4 = (K4rx84 | J1qx84);
	assign K4rx84 = (O9e2a4 & V9e2a4);
	assign V9e2a4 = (Cae2a4 & Jae2a4);
	assign Jae2a4 = (Qae2a4 & Xae2a4);
	assign Qae2a4 = (~(O3ux84 & Ebe2a4));
	assign Ebe2a4 = (~(Lbe2a4 & Sbe2a4));
	assign Sbe2a4 = (~(Zbe2a4 & R673a4[3]));
	assign Lbe2a4 = (~(Gce2a4 & K873a4[3]));
	assign Cae2a4 = (Nce2a4 & Uce2a4);
	assign Uce2a4 = (Ertx84 | Vkyx84);
	assign Nce2a4 = (Bde2a4 | Tjyx84);
	assign O9e2a4 = (Ide2a4 & Pde2a4);
	assign Pde2a4 = (Wde2a4 & Dee2a4);
	assign Dee2a4 = (~(Pu63a4[3] & Pttx84));
	assign Wde2a4 = (~(X473a4[3] & Yutx84));
	assign Ide2a4 = (Kee2a4 & Ree2a4);
	assign Ree2a4 = (~(HRDATA[3] & Fvtx84));
	assign Kee2a4 = (~(STCALIB[3] & Hwtx84));
	assign A9e2a4 = (Yee2a4 & Ffe2a4);
	assign Ffe2a4 = (M5rx84 | H0qx84);
	assign M5rx84 = (Mfe2a4 & Tfe2a4);
	assign Tfe2a4 = (Age2a4 & Hge2a4);
	assign Age2a4 = (~(Oge2a4 & Vge2a4));
	assign Mfe2a4 = (Che2a4 & Jhe2a4);
	assign Jhe2a4 = (~(Nnyx84 & V3ux84));
	assign Nnyx84 = (~(Qhe2a4 | Oge2a4));
	assign Qhe2a4 = (F5yx84 ? Eie2a4 : Xhe2a4);
	assign Che2a4 = (~(HRDATA[27] & Fvtx84));
	assign Yee2a4 = (R4rx84 | Rypx84);
	assign R4rx84 = (Lie2a4 & Sie2a4);
	assign Sie2a4 = (Zie2a4 & Gje2a4);
	assign Gje2a4 = (~(Pu63a4[11] & Pttx84));
	assign Zie2a4 = (Nje2a4 & Uje2a4);
	assign Uje2a4 = (Ertx84 | Tcyx84);
	assign Nje2a4 = (~(Bttx84 & Kbyx84));
	assign Lie2a4 = (Bke2a4 & Ike2a4);
	assign Ike2a4 = (~(STCALIB[11] & Hwtx84));
	assign Bke2a4 = (Pke2a4 & Wke2a4);
	assign Wke2a4 = (~(X473a4[11] & Yutx84));
	assign Pke2a4 = (~(HRDATA[11] & Fvtx84));
	assign M8e2a4 = (V0qx84 & Dle2a4);
	assign Dle2a4 = (T5rx84 | Tzpx84);
	assign T5rx84 = (Kle2a4 & Rle2a4);
	assign Rle2a4 = (Yle2a4 & Fme2a4);
	assign Fme2a4 = (Mme2a4 & Zrtx84);
	assign Mme2a4 = (~(Tme2a4 & Q7yx84));
	assign Yle2a4 = (Ane2a4 & Hne2a4);
	assign Hne2a4 = (Bde2a4 | H6yx84);
	assign Ane2a4 = (~(Pu63a4[19] & Pttx84));
	assign Kle2a4 = (One2a4 & Vne2a4);
	assign Vne2a4 = (~(STCALIB[19] & Hwtx84));
	assign One2a4 = (Coe2a4 & Joe2a4);
	assign Joe2a4 = (~(X473a4[19] & Yutx84));
	assign Coe2a4 = (~(HRDATA[19] & Fvtx84));
	assign R7e2a4 = (~(Qoe2a4 & Jq0x84));
	assign Gcax84 = (~(Xoe2a4 & Epe2a4));
	assign Epe2a4 = (~(Nj63a4[5] & Lpe2a4));
	assign Xoe2a4 = (Spe2a4 & Zpe2a4);
	assign Zpe2a4 = (F8e2a4 | U2kx84);
	assign U2kx84 = (Gqe2a4 & Nqe2a4);
	assign Nqe2a4 = (Uqe2a4 & Bre2a4);
	assign Bre2a4 = (Odrx84 | J1qx84);
	assign Odrx84 = (Ire2a4 & Pre2a4);
	assign Pre2a4 = (Wre2a4 & Dse2a4);
	assign Dse2a4 = (~(Pu63a4[5] & Pttx84));
	assign Wre2a4 = (Kse2a4 & Rse2a4);
	assign Rse2a4 = (Bde2a4 | Adyx84);
	assign Kse2a4 = (Ertx84 | Diyx84);
	assign Ire2a4 = (Yse2a4 & Fte2a4);
	assign Fte2a4 = (~(STCALIB[5] & Hwtx84));
	assign Yse2a4 = (Mte2a4 & Tte2a4);
	assign Tte2a4 = (~(X473a4[5] & Yutx84));
	assign Mte2a4 = (~(HRDATA[5] & Fvtx84));
	assign Uqe2a4 = (Aue2a4 & Hue2a4);
	assign Hue2a4 = (Qerx84 | H0qx84);
	assign Qerx84 = (Oue2a4 & Vue2a4);
	assign Vue2a4 = (~(HRDATA[29] & Fvtx84));
	assign Oue2a4 = (Cve2a4 & Hge2a4);
	assign Cve2a4 = (Jve2a4 | Vryx84);
	assign Vryx84 = (Qve2a4 & Xve2a4);
	assign Xve2a4 = (Ewe2a4 | Lwe2a4);
	assign Lwe2a4 = (Gxe2a4 ? Zwe2a4 : Swe2a4);
	assign Swe2a4 = (!Clyx84);
	assign Qve2a4 = (~(Woyx84 & Ewe2a4));
	assign Ewe2a4 = (Nxe2a4 | Uxe2a4);
	assign Uxe2a4 = (Bye2a4 & Iye2a4);
	assign Nxe2a4 = (~(Pye2a4 | Bye2a4));
	assign Aue2a4 = (Vdrx84 | Rypx84);
	assign Vdrx84 = (Wye2a4 & Dze2a4);
	assign Dze2a4 = (Kze2a4 & Rze2a4);
	assign Rze2a4 = (Yze2a4 & F0f2a4);
	assign F0f2a4 = (~(Gstx84 & Pijx84));
	assign Pijx84 = (~(M0f2a4 & T0f2a4));
	assign T0f2a4 = (A1f2a4 & H1f2a4);
	assign M0f2a4 = (O1f2a4 & R9c2a4);
	assign O1f2a4 = (Bgb2a4 | V1f2a4);
	assign Yze2a4 = (Ertx84 | Bayx84);
	assign Kze2a4 = (C2f2a4 & J2f2a4);
	assign J2f2a4 = (~(Bttx84 & Rbyx84));
	assign C2f2a4 = (~(Pu63a4[13] & Pttx84));
	assign Wye2a4 = (Q2f2a4 & X2f2a4);
	assign X2f2a4 = (~(STCALIB[13] & Hwtx84));
	assign Q2f2a4 = (E3f2a4 & L3f2a4);
	assign L3f2a4 = (~(X473a4[13] & Yutx84));
	assign E3f2a4 = (~(HRDATA[13] & Fvtx84));
	assign Gqe2a4 = (V0qx84 & S3f2a4);
	assign S3f2a4 = (Xerx84 | Tzpx84);
	assign Xerx84 = (Z3f2a4 & G4f2a4);
	assign G4f2a4 = (N4f2a4 & U4f2a4);
	assign U4f2a4 = (~(Pu63a4[21] & Pttx84));
	assign N4f2a4 = (B5f2a4 & I5f2a4);
	assign I5f2a4 = (Bde2a4 | A6yx84);
	assign B5f2a4 = (Ertx84 | K4yx84);
	assign Z3f2a4 = (P5f2a4 & W5f2a4);
	assign W5f2a4 = (~(STCALIB[21] & Hwtx84));
	assign P5f2a4 = (D6f2a4 & K6f2a4);
	assign K6f2a4 = (~(X473a4[21] & Yutx84));
	assign D6f2a4 = (~(HRDATA[21] & Fvtx84));
	assign Spe2a4 = (~(Qoe2a4 & Zt0x84));
	assign Zbax84 = (~(R6f2a4 & Y6f2a4));
	assign Y6f2a4 = (Tbb2a4 | Nocx84);
	assign R6f2a4 = (F7f2a4 & M7f2a4);
	assign M7f2a4 = (F8e2a4 | A5ex84);
	assign A5ex84 = (T7f2a4 & A8f2a4);
	assign A8f2a4 = (H8f2a4 & O8f2a4);
	assign O8f2a4 = (Noqx84 | J1qx84);
	assign Noqx84 = (V8f2a4 & C9f2a4);
	assign C9f2a4 = (J9f2a4 & Q9f2a4);
	assign Q9f2a4 = (~(Pu63a4[0] & Pttx84));
	assign J9f2a4 = (X9f2a4 & Eaf2a4);
	assign Eaf2a4 = (~(O3ux84 & Laf2a4));
	assign Laf2a4 = (~(Saf2a4 & Zaf2a4));
	assign Zaf2a4 = (~(Gce2a4 & K873a4[0]));
	assign Saf2a4 = (Gbf2a4 & Nbf2a4);
	assign Nbf2a4 = (~(Mq3x84 & W6hx84));
	assign Gbf2a4 = (~(Zbe2a4 & R673a4[0]));
	assign X9f2a4 = (~(Rqxx84 & V3ux84));
	assign Rqxx84 = (F5yx84 ? Bcf2a4 : Ubf2a4);
	assign V8f2a4 = (Icf2a4 & Pcf2a4);
	assign Pcf2a4 = (~(STCALIB[0] & Hwtx84));
	assign Icf2a4 = (Wcf2a4 & Ddf2a4);
	assign Ddf2a4 = (~(X473a4[0] & Yutx84));
	assign Wcf2a4 = (~(HRDATA[0] & Fvtx84));
	assign H8f2a4 = (Kdf2a4 & Rdf2a4);
	assign Rdf2a4 = (Dqqx84 | H0qx84);
	assign Dqqx84 = (Ydf2a4 & Fef2a4);
	assign Fef2a4 = (~(HRDATA[24] & Fvtx84));
	assign Ydf2a4 = (Mef2a4 & Zrtx84);
	assign Mef2a4 = (~(Unyx84 & V3ux84));
	assign Unyx84 = (Hsxx84 & Tef2a4);
	assign Tef2a4 = (Aff2a4 | Wlnx84);
	assign Hsxx84 = (Gxe2a4 ? O6yx84 : Hff2a4);
	assign Kdf2a4 = (Bpqx84 | Rypx84);
	assign Bpqx84 = (Off2a4 & Vff2a4);
	assign Vff2a4 = (Cgf2a4 & Jgf2a4);
	assign Jgf2a4 = (~(X473a4[8] & Yutx84));
	assign Cgf2a4 = (Qgf2a4 & Xgf2a4);
	assign Xgf2a4 = (~(Vsxx84 & V3ux84));
	assign Vsxx84 = (F5yx84 ? Mcyx84 : Mjyx84);
	assign Qgf2a4 = (~(Pu63a4[8] & Pttx84));
	assign Off2a4 = (Ehf2a4 & Lhf2a4);
	assign Lhf2a4 = (~(HRDATA[8] & Fvtx84));
	assign Ehf2a4 = (~(STCALIB[8] & Hwtx84));
	assign T7f2a4 = (V0qx84 & Shf2a4);
	assign Shf2a4 = (Rqqx84 | Tzpx84);
	assign Rqqx84 = (Zhf2a4 & Gif2a4);
	assign Gif2a4 = (Nif2a4 & Uif2a4);
	assign Uif2a4 = (Bjf2a4 & Hge2a4);
	assign Bjf2a4 = (~(Ijf2a4 & Vk3x84));
	assign Ijf2a4 = (W6hx84 & O3ux84);
	assign Nif2a4 = (Pjf2a4 & Wjf2a4);
	assign Wjf2a4 = (~(Aljx84 & Gstx84));
	assign Aljx84 = (Dkf2a4 & Ufb2a4);
	assign Pjf2a4 = (~(Asxx84 & V3ux84));
	assign Asxx84 = (F5yx84 ? J7yx84 : Dbyx84);
	assign Zhf2a4 = (Kkf2a4 & Rkf2a4);
	assign Rkf2a4 = (Ykf2a4 & Flf2a4);
	assign Flf2a4 = (~(Pu63a4[16] & Pttx84));
	assign Ykf2a4 = (~(X473a4[16] & Yutx84));
	assign Kkf2a4 = (Mlf2a4 & Tlf2a4);
	assign Tlf2a4 = (~(HRDATA[16] & Fvtx84));
	assign Mlf2a4 = (~(STCALIB[16] & Hwtx84));
	assign F7f2a4 = (~(Qoe2a4 & Yk0x84));
	assign Sbax84 = (~(Amf2a4 & Hmf2a4));
	assign Hmf2a4 = (Omf2a4 | Nocx84);
	assign Amf2a4 = (Vmf2a4 & Cnf2a4);
	assign Cnf2a4 = (F8e2a4 | Gygx84);
	assign Gygx84 = (Jnf2a4 & Qnf2a4);
	assign Qnf2a4 = (Xnf2a4 & Eof2a4);
	assign Eof2a4 = (J1qx84 | Qtqx84);
	assign Qtqx84 = (Lof2a4 & Sof2a4);
	assign Sof2a4 = (Zof2a4 & Gpf2a4);
	assign Gpf2a4 = (Npf2a4 & Upf2a4);
	assign Upf2a4 = (~(O3ux84 & Bqf2a4));
	assign Bqf2a4 = (~(Iqf2a4 & Pqf2a4));
	assign Pqf2a4 = (Wqf2a4 & Drf2a4);
	assign Drf2a4 = (~(Krf2a4 & M8hx84));
	assign Krf2a4 = (V2hx84 & Lo4w84);
	assign Wqf2a4 = (~(Oo3x84 & W6hx84));
	assign Iqf2a4 = (Rrf2a4 & Yrf2a4);
	assign Yrf2a4 = (~(Zbe2a4 & R673a4[1]));
	assign Rrf2a4 = (~(Gce2a4 & K873a4[1]));
	assign Npf2a4 = (~(Tme2a4 & Clyx84));
	assign Clyx84 = (~(Fsf2a4 & Msf2a4));
	assign Msf2a4 = (Tsf2a4 & Atf2a4);
	assign Atf2a4 = (~(Htf2a4 & Otf2a4));
	assign Tsf2a4 = (~(Aryx84 & Vtf2a4));
	assign Fsf2a4 = (Cuf2a4 & Juf2a4);
	assign Juf2a4 = (~(Quf2a4 & Xuf2a4));
	assign Cuf2a4 = (~(Tqyx84 & Evf2a4));
	assign Zof2a4 = (Lvf2a4 & Svf2a4);
	assign Svf2a4 = (Bde2a4 | Diyx84);
	assign Diyx84 = (Zvf2a4 & Gwf2a4);
	assign Gwf2a4 = (Nwf2a4 & Uwf2a4);
	assign Uwf2a4 = (~(Htf2a4 & Bxf2a4));
	assign Nwf2a4 = (~(Aryx84 & Ixf2a4));
	assign Zvf2a4 = (Pxf2a4 & Wxf2a4);
	assign Wxf2a4 = (~(Quf2a4 & Dyf2a4));
	assign Pxf2a4 = (~(Tqyx84 & Kyf2a4));
	assign Lvf2a4 = (~(Pu63a4[1] & Pttx84));
	assign Lof2a4 = (Ryf2a4 & Yyf2a4);
	assign Yyf2a4 = (~(STCALIB[1] & Hwtx84));
	assign Ryf2a4 = (Fzf2a4 & Mzf2a4);
	assign Mzf2a4 = (~(X473a4[1] & Yutx84));
	assign Fzf2a4 = (~(HRDATA[1] & Fvtx84));
	assign Xnf2a4 = (Tzf2a4 & A0g2a4);
	assign A0g2a4 = (H0qx84 | Luqx84);
	assign Luqx84 = (H0g2a4 & O0g2a4);
	assign O0g2a4 = (V0g2a4 & Hge2a4);
	assign V0g2a4 = (~(Vge2a4 & C1g2a4));
	assign H0g2a4 = (J1g2a4 & Q1g2a4);
	assign Q1g2a4 = (~(Gnyx84 & V3ux84));
	assign Gnyx84 = (~(X1g2a4 | C1g2a4));
	assign C1g2a4 = (E2g2a4 & L2g2a4);
	assign E2g2a4 = (Aff2a4 ? Bye2a4 : S2g2a4);
	assign S2g2a4 = (~(Z2g2a4 & Bye2a4));
	assign Bye2a4 = (~(Quf2a4 | Aryx84));
	assign X1g2a4 = (F5yx84 ? Zwe2a4 : A6yx84);
	assign Zwe2a4 = (G3g2a4 & N3g2a4);
	assign N3g2a4 = (U3g2a4 & B4g2a4);
	assign B4g2a4 = (~(Htf2a4 & I4g2a4));
	assign U3g2a4 = (~(Aryx84 & P4g2a4));
	assign G3g2a4 = (W4g2a4 & D5g2a4);
	assign D5g2a4 = (~(Quf2a4 & K5g2a4));
	assign W4g2a4 = (~(Tqyx84 & R5g2a4));
	assign A6yx84 = (Y5g2a4 & F6g2a4);
	assign F6g2a4 = (M6g2a4 & T6g2a4);
	assign T6g2a4 = (~(Htf2a4 & A7g2a4));
	assign M6g2a4 = (~(Aryx84 & H7g2a4));
	assign Y5g2a4 = (O7g2a4 & V7g2a4);
	assign V7g2a4 = (~(Quf2a4 & C8g2a4));
	assign O7g2a4 = (~(Tqyx84 & J8g2a4));
	assign J1g2a4 = (~(HRDATA[25] & Fvtx84));
	assign Tzf2a4 = (Rypx84 | Ctqx84);
	assign Ctqx84 = (Q8g2a4 & X8g2a4);
	assign X8g2a4 = (E9g2a4 & L9g2a4);
	assign L9g2a4 = (Zrtx84 & Xae2a4);
	assign Xae2a4 = (~(S9g2a4 & Z9g2a4));
	assign E9g2a4 = (Gag2a4 & Nag2a4);
	assign Nag2a4 = (Ertx84 | Adyx84);
	assign Adyx84 = (Uag2a4 & Bbg2a4);
	assign Bbg2a4 = (Ibg2a4 & Pbg2a4);
	assign Pbg2a4 = (~(Htf2a4 & Wbg2a4));
	assign Ibg2a4 = (~(Aryx84 & Dcg2a4));
	assign Uag2a4 = (Kcg2a4 & Rcg2a4);
	assign Rcg2a4 = (~(Quf2a4 & Ycg2a4));
	assign Kcg2a4 = (~(Tqyx84 & Fdg2a4));
	assign Ertx84 = (!Tme2a4);
	assign Gag2a4 = (Bde2a4 | Bayx84);
	assign Bayx84 = (Mdg2a4 & Tdg2a4);
	assign Tdg2a4 = (Aeg2a4 & Heg2a4);
	assign Heg2a4 = (~(Htf2a4 & Oeg2a4));
	assign Aeg2a4 = (~(Aryx84 & Veg2a4));
	assign Mdg2a4 = (Cfg2a4 & Jfg2a4);
	assign Jfg2a4 = (~(Quf2a4 & Qfg2a4));
	assign Cfg2a4 = (~(Tqyx84 & Xfg2a4));
	assign Q8g2a4 = (Egg2a4 & Lgg2a4);
	assign Lgg2a4 = (Sgg2a4 & Zgg2a4);
	assign Zgg2a4 = (~(Pu63a4[9] & Pttx84));
	assign Sgg2a4 = (~(X473a4[9] & Yutx84));
	assign Egg2a4 = (Ghg2a4 & Nhg2a4);
	assign Nhg2a4 = (~(HRDATA[9] & Fvtx84));
	assign Ghg2a4 = (~(STCALIB[9] & Hwtx84));
	assign Jnf2a4 = (V0qx84 & Uhg2a4);
	assign Uhg2a4 = (Tzpx84 | Suqx84);
	assign Suqx84 = (Big2a4 & Iig2a4);
	assign Iig2a4 = (Pig2a4 & Wig2a4);
	assign Wig2a4 = (~(Pu63a4[17] & Pttx84));
	assign Pig2a4 = (Djg2a4 & Kjg2a4);
	assign Kjg2a4 = (~(Tme2a4 & Rbyx84));
	assign Rbyx84 = (~(Rjg2a4 & Yjg2a4));
	assign Yjg2a4 = (Fkg2a4 & Mkg2a4);
	assign Mkg2a4 = (~(Htf2a4 & Tkg2a4));
	assign Fkg2a4 = (~(Aryx84 & Alg2a4));
	assign Rjg2a4 = (Hlg2a4 & Olg2a4);
	assign Olg2a4 = (~(Quf2a4 & Vlg2a4));
	assign Hlg2a4 = (~(Tqyx84 & Cmg2a4));
	assign Djg2a4 = (Bde2a4 | K4yx84);
	assign K4yx84 = (Jmg2a4 & Qmg2a4);
	assign Qmg2a4 = (Xmg2a4 & Eng2a4);
	assign Eng2a4 = (~(Htf2a4 & Lng2a4));
	assign Xmg2a4 = (~(Aryx84 & Sng2a4));
	assign Jmg2a4 = (Zng2a4 & Gog2a4);
	assign Gog2a4 = (~(Quf2a4 & Nog2a4));
	assign Zng2a4 = (~(Tqyx84 & Uog2a4));
	assign Big2a4 = (Bpg2a4 & Ipg2a4);
	assign Ipg2a4 = (~(STCALIB[17] & Hwtx84));
	assign Bpg2a4 = (Ppg2a4 & Wpg2a4);
	assign Wpg2a4 = (~(X473a4[17] & Yutx84));
	assign Ppg2a4 = (~(HRDATA[17] & Fvtx84));
	assign Vmf2a4 = (~(Qoe2a4 & Tm0x84));
	assign Lbax84 = (~(Dqg2a4 & Kqg2a4));
	assign Kqg2a4 = (Rqg2a4 | Nocx84);
	assign Dqg2a4 = (Yqg2a4 & Frg2a4);
	assign Frg2a4 = (F8e2a4 | G9kx84);
	assign G9kx84 = (Mrg2a4 & Trg2a4);
	assign Trg2a4 = (Asg2a4 & Hsg2a4);
	assign Hsg2a4 = (Hzqx84 | J1qx84);
	assign Hzqx84 = (Osg2a4 & Vsg2a4);
	assign Vsg2a4 = (Ctg2a4 & Jtg2a4);
	assign Jtg2a4 = (Qtg2a4 & Xtg2a4);
	assign Xtg2a4 = (~(O3ux84 & Eug2a4));
	assign Eug2a4 = (~(Lug2a4 & Sug2a4));
	assign Sug2a4 = (Zug2a4 & Gvg2a4);
	assign Gvg2a4 = (~(Nvg2a4 & Y63x84));
	assign Nvg2a4 = (M8hx84 & V2hx84);
	assign Zug2a4 = (~(W6hx84 & P6e2a4));
	assign P6e2a4 = (Qm3x84 | STCALIB[25]);
	assign W6hx84 = (R7hx84 & J0kx84);
	assign Lug2a4 = (Uvg2a4 & Bwg2a4);
	assign Bwg2a4 = (~(Zbe2a4 & R673a4[2]));
	assign Zbe2a4 = (I6hx84 & Iwg2a4);
	assign Uvg2a4 = (~(Gce2a4 & K873a4[2]));
	assign Gce2a4 = (T8hx84 & Iwg2a4);
	assign Iwg2a4 = (J0kx84 | Fhfx84);
	assign Qtg2a4 = (~(Tme2a4 & Jlyx84));
	assign Jlyx84 = (~(Pwg2a4 & Wwg2a4));
	assign Wwg2a4 = (Dxg2a4 & Kxg2a4);
	assign Kxg2a4 = (~(Htf2a4 & Kyf2a4));
	assign Dxg2a4 = (~(Aryx84 & Xuf2a4));
	assign Pwg2a4 = (Rxg2a4 & Yxg2a4);
	assign Yxg2a4 = (~(Quf2a4 & Otf2a4));
	assign Rxg2a4 = (~(Tqyx84 & Vtf2a4));
	assign Ctg2a4 = (Fyg2a4 & Myg2a4);
	assign Myg2a4 = (Bde2a4 | D8ux84);
	assign D8ux84 = (Tyg2a4 & Azg2a4);
	assign Azg2a4 = (Hzg2a4 & Ozg2a4);
	assign Ozg2a4 = (~(Htf2a4 & Fdg2a4));
	assign Hzg2a4 = (~(Aryx84 & Dyf2a4));
	assign Tyg2a4 = (Vzg2a4 & C0h2a4);
	assign C0h2a4 = (~(Quf2a4 & Bxf2a4));
	assign Vzg2a4 = (~(Tqyx84 & Ixf2a4));
	assign Fyg2a4 = (~(Pu63a4[2] & Pttx84));
	assign Osg2a4 = (J0h2a4 & Q0h2a4);
	assign Q0h2a4 = (~(STCALIB[2] & Hwtx84));
	assign J0h2a4 = (X0h2a4 & E1h2a4);
	assign E1h2a4 = (~(X473a4[2] & Yutx84));
	assign X0h2a4 = (~(HRDATA[2] & Fvtx84));
	assign Asg2a4 = (L1h2a4 & S1h2a4);
	assign S1h2a4 = (J0rx84 | H0qx84);
	assign J0rx84 = (Z1h2a4 & G2h2a4);
	assign G2h2a4 = (~(HRDATA[26] & Fvtx84));
	assign Z1h2a4 = (N2h2a4 & U2h2a4);
	assign U2h2a4 = (Jve2a4 | Csyx84);
	assign Csyx84 = (B3h2a4 & I3h2a4);
	assign I3h2a4 = (~(Oge2a4 & Woyx84));
	assign B3h2a4 = (P3h2a4 | W3h2a4);
	assign W3h2a4 = (Aryx84 ? D4h2a4 : Oge2a4);
	assign D4h2a4 = (L2g2a4 & K4h2a4);
	assign Oge2a4 = (L2g2a4 & R4h2a4);
	assign R4h2a4 = (~(Z2g2a4 & K4h2a4));
	assign L2g2a4 = (Y4h2a4 & Wbcx84);
	assign Y4h2a4 = (K4h2a4 | Z2g2a4);
	assign Z2g2a4 = (F5yx84 & F5h2a4);
	assign P3h2a4 = (!M5h2a4);
	assign M5h2a4 = (Gxe2a4 ? Sytx84 : Oryx84);
	assign Sytx84 = (~(T5h2a4 & A6h2a4));
	assign A6h2a4 = (H6h2a4 & O6h2a4);
	assign O6h2a4 = (~(Htf2a4 & R5g2a4));
	assign H6h2a4 = (~(Aryx84 & C8g2a4));
	assign T5h2a4 = (V6h2a4 & C7h2a4);
	assign C7h2a4 = (~(Quf2a4 & A7g2a4));
	assign V6h2a4 = (~(Tqyx84 & H7g2a4));
	assign Oryx84 = (~(J7h2a4 & Q7h2a4));
	assign Q7h2a4 = (X7h2a4 & E8h2a4);
	assign E8h2a4 = (~(Htf2a4 & Evf2a4));
	assign X7h2a4 = (~(Aryx84 & K5g2a4));
	assign J7h2a4 = (L8h2a4 & S8h2a4);
	assign S8h2a4 = (~(Quf2a4 & I4g2a4));
	assign L8h2a4 = (~(Tqyx84 & P4g2a4));
	assign N2h2a4 = (~(Gstx84 & Js3x84));
	assign L1h2a4 = (Ozqx84 | Rypx84);
	assign Ozqx84 = (Z8h2a4 & G9h2a4);
	assign G9h2a4 = (N9h2a4 & U9h2a4);
	assign U9h2a4 = (~(Pu63a4[10] & Pttx84));
	assign N9h2a4 = (Bah2a4 & Iah2a4);
	assign Iah2a4 = (~(Tme2a4 & W7ux84));
	assign W7ux84 = (~(Pah2a4 & Wah2a4));
	assign Wah2a4 = (Dbh2a4 & Kbh2a4);
	assign Kbh2a4 = (~(Htf2a4 & Xfg2a4));
	assign Dbh2a4 = (~(Aryx84 & Ycg2a4));
	assign Pah2a4 = (Rbh2a4 & Ybh2a4);
	assign Ybh2a4 = (~(Quf2a4 & Wbg2a4));
	assign Rbh2a4 = (~(Tqyx84 & Dcg2a4));
	assign Bah2a4 = (Bde2a4 | Lrtx84);
	assign Lrtx84 = (Fch2a4 & Mch2a4);
	assign Mch2a4 = (Tch2a4 & Adh2a4);
	assign Adh2a4 = (~(Htf2a4 & Cmg2a4));
	assign Tch2a4 = (~(Aryx84 & Qfg2a4));
	assign Fch2a4 = (Hdh2a4 & Odh2a4);
	assign Odh2a4 = (~(Quf2a4 & Oeg2a4));
	assign Hdh2a4 = (~(Tqyx84 & Veg2a4));
	assign Z8h2a4 = (Vdh2a4 & Ceh2a4);
	assign Ceh2a4 = (~(STCALIB[10] & Hwtx84));
	assign Vdh2a4 = (Jeh2a4 & Qeh2a4);
	assign Qeh2a4 = (~(X473a4[10] & Yutx84));
	assign Jeh2a4 = (~(HRDATA[10] & Fvtx84));
	assign Mrg2a4 = (V0qx84 & Xeh2a4);
	assign Xeh2a4 = (Q0rx84 | Tzpx84);
	assign Q0rx84 = (Efh2a4 & Lfh2a4);
	assign Lfh2a4 = (Sfh2a4 & M2ux84);
	assign M2ux84 = (Hge2a4 & Zrtx84);
	assign Sfh2a4 = (Zfh2a4 & Ggh2a4);
	assign Ggh2a4 = (~(Tme2a4 & Ittx84));
	assign Ittx84 = (~(Ngh2a4 & Ugh2a4));
	assign Ugh2a4 = (Bhh2a4 & Ihh2a4);
	assign Ihh2a4 = (~(Htf2a4 & Uog2a4));
	assign Bhh2a4 = (~(Aryx84 & Vlg2a4));
	assign Ngh2a4 = (Phh2a4 & Whh2a4);
	assign Whh2a4 = (~(Quf2a4 & Tkg2a4));
	assign Phh2a4 = (~(Tqyx84 & Alg2a4));
	assign Zfh2a4 = (Bde2a4 | Zytx84);
	assign Zytx84 = (Dih2a4 & Kih2a4);
	assign Kih2a4 = (Rih2a4 & Yih2a4);
	assign Yih2a4 = (~(Htf2a4 & J8g2a4));
	assign Rih2a4 = (~(Aryx84 & Nog2a4));
	assign Dih2a4 = (Fjh2a4 & Mjh2a4);
	assign Mjh2a4 = (~(Quf2a4 & Lng2a4));
	assign Fjh2a4 = (~(Tqyx84 & Sng2a4));
	assign Bde2a4 = (!Bttx84);
	assign Efh2a4 = (Tjh2a4 & Akh2a4);
	assign Akh2a4 = (Hkh2a4 & Okh2a4);
	assign Okh2a4 = (~(Pu63a4[18] & Pttx84));
	assign Hkh2a4 = (~(X473a4[18] & Yutx84));
	assign Tjh2a4 = (Vkh2a4 & Clh2a4);
	assign Clh2a4 = (~(HRDATA[18] & Fvtx84));
	assign Vkh2a4 = (~(STCALIB[18] & Hwtx84));
	assign Yqg2a4 = (~(Qoe2a4 & Oo0x84));
	assign Ebax84 = (~(Jlh2a4 & Qlh2a4));
	assign Qlh2a4 = (~(Nj63a4[4] & Lpe2a4));
	assign Lpe2a4 = (!Nocx84);
	assign Jlh2a4 = (Xlh2a4 & Emh2a4);
	assign Emh2a4 = (F8e2a4 | O7qx84);
	assign O7qx84 = (Lmh2a4 & Smh2a4);
	assign Smh2a4 = (Zmh2a4 & Gnh2a4);
	assign Gnh2a4 = (E8rx84 | J1qx84);
	assign J1qx84 = (Iorx84 & Nnh2a4);
	assign Nnh2a4 = (~(Unh2a4 & Orrx84));
	assign Unh2a4 = (~(Boh2a4 & Ioh2a4));
	assign Ioh2a4 = (M6xx84 | Zo2x84);
	assign Boh2a4 = (Poh2a4 & Woh2a4);
	assign Woh2a4 = (~(Dph2a4 & Kph2a4));
	assign Kph2a4 = (Ns2x84 | Mbex84);
	assign Poh2a4 = (W1c2a4 | Kshx84);
	assign Iorx84 = (Hhux84 | Rph2a4);
	assign Rph2a4 = (Yph2a4 & Fqh2a4);
	assign Fqh2a4 = (~(Rprx84 | Uwix84));
	assign Yph2a4 = (~(Gpbx84 | Tsix84));
	assign E8rx84 = (Mqh2a4 & Tqh2a4);
	assign Tqh2a4 = (Arh2a4 & Hrh2a4);
	assign Hrh2a4 = (Orh2a4 & Vrh2a4);
	assign Vrh2a4 = (~(Csh2a4 & R83x84));
	assign Csh2a4 = (M8hx84 & S9g2a4);
	assign Orh2a4 = (~(Tme2a4 & Bcf2a4));
	assign Bcf2a4 = (!Okyx84);
	assign Okyx84 = (Jsh2a4 & Qsh2a4);
	assign Qsh2a4 = (Xsh2a4 & Eth2a4);
	assign Eth2a4 = (~(Htf2a4 & Dyf2a4));
	assign Xsh2a4 = (~(Aryx84 & Kyf2a4));
	assign Jsh2a4 = (Lth2a4 & Sth2a4);
	assign Sth2a4 = (~(Quf2a4 & Ixf2a4));
	assign Lth2a4 = (~(Tqyx84 & Otf2a4));
	assign Arh2a4 = (Zth2a4 & Guh2a4);
	assign Guh2a4 = (~(Bttx84 & Mjyx84));
	assign Mjyx84 = (~(Nuh2a4 & Uuh2a4));
	assign Uuh2a4 = (Bvh2a4 & Ivh2a4);
	assign Ivh2a4 = (~(Htf2a4 & Ycg2a4));
	assign Bvh2a4 = (~(Quf2a4 & Dcg2a4));
	assign Nuh2a4 = (Pvh2a4 & Wvh2a4);
	assign Wvh2a4 = (~(Aryx84 & Fdg2a4));
	assign Pvh2a4 = (~(Tqyx84 & Bxf2a4));
	assign Zth2a4 = (~(Pu63a4[4] & Pttx84));
	assign Mqh2a4 = (Dwh2a4 & Kwh2a4);
	assign Kwh2a4 = (~(STCALIB[4] & Hwtx84));
	assign Dwh2a4 = (Rwh2a4 & Ywh2a4);
	assign Ywh2a4 = (~(X473a4[4] & Yutx84));
	assign Rwh2a4 = (~(HRDATA[4] & Fvtx84));
	assign Zmh2a4 = (Fxh2a4 & Mxh2a4);
	assign Mxh2a4 = (G9rx84 | H0qx84);
	assign H0qx84 = (Txh2a4 & Ayh2a4);
	assign Ayh2a4 = (~(Hyh2a4 & Vs63a4[1]));
	assign Txh2a4 = (Oyh2a4 & Qsrx84);
	assign Qsrx84 = (F5dx84 | Rprx84);
	assign Oyh2a4 = (Sfyx84 | Orrx84);
	assign G9rx84 = (Vyh2a4 & Czh2a4);
	assign Czh2a4 = (Jzh2a4 & Hge2a4);
	assign Jzh2a4 = (~(V3ux84 & Poyx84));
	assign Poyx84 = (Pye2a4 ? Qzh2a4 : Woyx84);
	assign Qzh2a4 = (F5yx84 ? Ubf2a4 : Hff2a4);
	assign Ubf2a4 = (~(Xzh2a4 & E0i2a4));
	assign E0i2a4 = (L0i2a4 & S0i2a4);
	assign S0i2a4 = (~(Htf2a4 & Xuf2a4));
	assign L0i2a4 = (~(Aryx84 & Evf2a4));
	assign Xzh2a4 = (Z0i2a4 & G1i2a4);
	assign G1i2a4 = (~(Quf2a4 & Vtf2a4));
	assign Z0i2a4 = (~(Tqyx84 & I4g2a4));
	assign Hff2a4 = (~(N1i2a4 & U1i2a4));
	assign U1i2a4 = (B2i2a4 & I2i2a4);
	assign I2i2a4 = (~(Htf2a4 & K5g2a4));
	assign B2i2a4 = (~(Aryx84 & R5g2a4));
	assign N1i2a4 = (P2i2a4 & W2i2a4);
	assign W2i2a4 = (~(Quf2a4 & P4g2a4));
	assign P2i2a4 = (~(Tqyx84 & A7g2a4));
	assign Vyh2a4 = (D3i2a4 & K3i2a4);
	assign K3i2a4 = (~(Gstx84 & Td3x84));
	assign D3i2a4 = (~(HRDATA[28] & Fvtx84));
	assign Fxh2a4 = (L8rx84 | Rypx84);
	assign Rypx84 = (R3i2a4 & Borx84);
	assign Borx84 = (~(Y3i2a4 & Orrx84));
	assign R3i2a4 = (F4i2a4 & Xsrx84);
	assign Xsrx84 = (Odyx84 | Orrx84);
	assign F4i2a4 = (~(Hyh2a4 & M4i2a4));
	assign M4i2a4 = (!Vs63a4[1]);
	assign Hyh2a4 = (T4i2a4 & Vs63a4[0]);
	assign T4i2a4 = (~(Xqfx84 | Rprx84));
	assign Xqfx84 = (Wqbx84 | J13x84);
	assign L8rx84 = (A5i2a4 & H5i2a4);
	assign H5i2a4 = (O5i2a4 & V5i2a4);
	assign V5i2a4 = (C6i2a4 & J6i2a4);
	assign J6i2a4 = (~(Yjjx84 & Gstx84));
	assign Yjjx84 = (Q6i2a4 & Mhfx84);
	assign Mhfx84 = (!La3x84);
	assign Q6i2a4 = (X6i2a4 | Cc3x84);
	assign X6i2a4 = (Pgb2a4 ? L7i2a4 : E7i2a4);
	assign E7i2a4 = (S7i2a4 & Nj72a4);
	assign S7i2a4 = (Z7i2a4 | Bgb2a4);
	assign Z7i2a4 = (V1f2a4 ? N8i2a4 : G8i2a4);
	assign C6i2a4 = (~(Tme2a4 & Mcyx84));
	assign Mcyx84 = (~(U8i2a4 & B9i2a4));
	assign B9i2a4 = (I9i2a4 & P9i2a4);
	assign P9i2a4 = (~(Quf2a4 & Veg2a4));
	assign I9i2a4 = (~(Htf2a4 & Qfg2a4));
	assign U8i2a4 = (W9i2a4 & Dai2a4);
	assign Dai2a4 = (~(Aryx84 & Xfg2a4));
	assign W9i2a4 = (~(Tqyx84 & Wbg2a4));
	assign O5i2a4 = (Kai2a4 & Rai2a4);
	assign Rai2a4 = (~(Bttx84 & Dbyx84));
	assign Dbyx84 = (~(Yai2a4 & Fbi2a4));
	assign Fbi2a4 = (Mbi2a4 & Tbi2a4);
	assign Tbi2a4 = (~(Htf2a4 & Vlg2a4));
	assign Mbi2a4 = (~(Aryx84 & Cmg2a4));
	assign Yai2a4 = (Aci2a4 & Hci2a4);
	assign Hci2a4 = (~(Quf2a4 & Alg2a4));
	assign Aci2a4 = (~(Tqyx84 & Oeg2a4));
	assign Kai2a4 = (~(Pu63a4[12] & Pttx84));
	assign A5i2a4 = (Oci2a4 & Vci2a4);
	assign Vci2a4 = (~(STCALIB[12] & Hwtx84));
	assign Oci2a4 = (Cdi2a4 & Jdi2a4);
	assign Jdi2a4 = (~(X473a4[12] & Yutx84));
	assign Cdi2a4 = (~(HRDATA[12] & Fvtx84));
	assign Lmh2a4 = (V0qx84 & Qdi2a4);
	assign Qdi2a4 = (N9rx84 | Tzpx84);
	assign Tzpx84 = (Xdi2a4 & Eei2a4);
	assign Eei2a4 = (~(Lei2a4 & Sei2a4));
	assign Sei2a4 = (Zei2a4 & Orrx84);
	assign Zei2a4 = (~(Vs63a4[0] | J13x84));
	assign Lei2a4 = (Vs63a4[1] & Gfi2a4);
	assign Gfi2a4 = (~(Wqbx84 & Nfi2a4));
	assign Nfi2a4 = (~(Zvix84 & Qxmx84));
	assign Xdi2a4 = (Mqrx84 | Ufi2a4);
	assign Mqrx84 = (Bgi2a4 | Orrx84);
	assign N9rx84 = (Igi2a4 & Pgi2a4);
	assign Pgi2a4 = (Wgi2a4 & Dhi2a4);
	assign Dhi2a4 = (~(Pu63a4[20] & Pttx84));
	assign Wgi2a4 = (Khi2a4 & Rhi2a4);
	assign Rhi2a4 = (~(Tme2a4 & J7yx84));
	assign J7yx84 = (~(Yhi2a4 & Fii2a4));
	assign Fii2a4 = (Mii2a4 & Tii2a4);
	assign Tii2a4 = (~(Htf2a4 & Nog2a4));
	assign Mii2a4 = (~(Aryx84 & Uog2a4));
	assign Yhi2a4 = (Aji2a4 & Hji2a4);
	assign Hji2a4 = (~(Quf2a4 & Sng2a4));
	assign Aji2a4 = (~(Tqyx84 & Tkg2a4));
	assign Tme2a4 = (~(Jve2a4 | F5yx84));
	assign Khi2a4 = (~(Bttx84 & O6yx84));
	assign O6yx84 = (~(Oji2a4 & Vji2a4));
	assign Vji2a4 = (Cki2a4 & Jki2a4);
	assign Jki2a4 = (~(Htf2a4 & C8g2a4));
	assign Cki2a4 = (~(Aryx84 & J8g2a4));
	assign Oji2a4 = (Qki2a4 & Xki2a4);
	assign Xki2a4 = (~(Quf2a4 & H7g2a4));
	assign Qki2a4 = (~(Tqyx84 & Lng2a4));
	assign Bttx84 = (~(Jve2a4 | Gxe2a4));
	assign Igi2a4 = (Eli2a4 & Lli2a4);
	assign Lli2a4 = (~(STCALIB[20] & Hwtx84));
	assign Eli2a4 = (Sli2a4 & Zli2a4);
	assign Zli2a4 = (~(X473a4[20] & Yutx84));
	assign Sli2a4 = (~(HRDATA[20] & Fvtx84));
	assign V0qx84 = (Gmi2a4 & Nmi2a4);
	assign Nmi2a4 = (~(Umi2a4 & Bni2a4));
	assign Bni2a4 = (X7yx84 & Sfyx84);
	assign Sfyx84 = (~(Ini2a4 & Olxx84));
	assign Ini2a4 = (~(Cmxx84 | Pni2a4));
	assign X7yx84 = (Wni2a4 & Odyx84);
	assign Odyx84 = (Fgux84 | Ufi2a4);
	assign Fgux84 = (~(Doi2a4 & Osxx84));
	assign Doi2a4 = (~(Pni2a4 | Olxx84));
	assign Wni2a4 = (Bgi2a4 | Ufi2a4);
	assign Bgi2a4 = (!Ngyx84);
	assign Ngyx84 = (Koi2a4 & Olxx84);
	assign Koi2a4 = (~(Pni2a4 | Osxx84));
	assign Pni2a4 = (!Xlyx84);
	assign Umi2a4 = (Hhux84 & Gurx84);
	assign Gurx84 = (~(Roi2a4 & Yoi2a4));
	assign Yoi2a4 = (Fpi2a4 & Mpi2a4);
	assign Mpi2a4 = (~(Tpi2a4 & Pz2x84));
	assign Tpi2a4 = (~(Aqi2a4 | Mkqx84));
	assign Mkqx84 = (Hqi2a4 & Oqi2a4);
	assign Oqi2a4 = (Vqi2a4 & Cri2a4);
	assign Cri2a4 = (~(X473a4[7] & Yutx84));
	assign Vqi2a4 = (Jri2a4 & Qri2a4);
	assign Qri2a4 = (Jve2a4 | Suxx84);
	assign Suxx84 = (F5yx84 ? Tcyx84 : Tjyx84);
	assign Tcyx84 = (Xri2a4 & Esi2a4);
	assign Esi2a4 = (Lsi2a4 & Ssi2a4);
	assign Ssi2a4 = (~(Quf2a4 & Xfg2a4));
	assign Lsi2a4 = (~(Tqyx84 & Ycg2a4));
	assign Xri2a4 = (Zsi2a4 & Gti2a4);
	assign Gti2a4 = (~(Htf2a4 & Veg2a4));
	assign Zsi2a4 = (~(Aryx84 & Wbg2a4));
	assign Tjyx84 = (Nti2a4 & Uti2a4);
	assign Uti2a4 = (Bui2a4 & Iui2a4);
	assign Iui2a4 = (~(Quf2a4 & Fdg2a4));
	assign Bui2a4 = (~(Tqyx84 & Dyf2a4));
	assign Nti2a4 = (Pui2a4 & Wui2a4);
	assign Wui2a4 = (~(Htf2a4 & Dcg2a4));
	assign Pui2a4 = (~(Aryx84 & Bxf2a4));
	assign Jri2a4 = (~(Pu63a4[7] & Pttx84));
	assign Hqi2a4 = (Dvi2a4 & Kvi2a4);
	assign Kvi2a4 = (~(STCALIB[7] & Hwtx84));
	assign Dvi2a4 = (Rvi2a4 & Yvi2a4);
	assign Yvi2a4 = (~(HRDATA[7] & Fvtx84));
	assign Rvi2a4 = (~(Nz63a4[1] & Awtx84));
	assign Aqi2a4 = (Fwi2a4 & Mwi2a4);
	assign Mwi2a4 = (~(Dph2a4 & Mgnx84));
	assign Dph2a4 = (~(Vs63a4[0] | Vs63a4[1]));
	assign Fwi2a4 = (Kshx84 | Qxmx84);
	assign Fpi2a4 = (Luxx84 & Pvrx84);
	assign Roi2a4 = (Twi2a4 & Axi2a4);
	assign Axi2a4 = (Hxi2a4 | Olqx84);
	assign Olqx84 = (Oxi2a4 & Vxi2a4);
	assign Vxi2a4 = (Cyi2a4 & Jyi2a4);
	assign Jyi2a4 = (Qyi2a4 & Zrtx84);
	assign Zrtx84 = (~(Xyi2a4 & M8hx84));
	assign Xyi2a4 = (O3ux84 & I6hx84);
	assign Qyi2a4 = (~(Gstx84 & Tkjx84));
	assign Tkjx84 = (~(Ezi2a4 | Dkf2a4));
	assign Dkf2a4 = (~(Bgb2a4 | Pgb2a4));
	assign Pgb2a4 = (!R9c2a4);
	assign Ezi2a4 = (!Ufb2a4);
	assign Ufb2a4 = (A1f2a4 & Nj72a4);
	assign Nj72a4 = (~(Lzi2a4 & R9c2a4));
	assign R9c2a4 = (~(Szi2a4 & Zzi2a4));
	assign Zzi2a4 = (L7i2a4 | Td3x84);
	assign Szi2a4 = (~(G0j2a4 & N0j2a4));
	assign N0j2a4 = (U0j2a4 & B1j2a4);
	assign B1j2a4 = (~(K9c2a4 & I1j2a4));
	assign I1j2a4 = (~(P1j2a4 & D9c2a4));
	assign P1j2a4 = (W1j2a4 & L6c2a4);
	assign L6c2a4 = (Igb2a4 ? Hw63a4[0] : Xx63a4[0]);
	assign K9c2a4 = (H1f2a4 ? D2j2a4 : D373a4[1]);
	assign U0j2a4 = (W1j2a4 | D9c2a4);
	assign D9c2a4 = (Igb2a4 ? Hw63a4[1] : Xx63a4[1]);
	assign W1j2a4 = (!E6c2a4);
	assign E6c2a4 = (H1f2a4 ? K2j2a4 : D373a4[0]);
	assign G0j2a4 = (R2j2a4 & Y2j2a4);
	assign Y2j2a4 = (~(H1f2a4 & Bgb2a4));
	assign R2j2a4 = (L7i2a4 ? M3j2a4 : F3j2a4);
	assign L7i2a4 = (!Igb2a4);
	assign Igb2a4 = (~(Kf3x84 & T3j2a4));
	assign T3j2a4 = (~(A4j2a4 & Td3x84));
	assign A4j2a4 = (H4j2a4 & O4j2a4);
	assign O4j2a4 = (Xx63a4[1] | V4j2a4);
	assign V4j2a4 = (C5j2a4 & Xx63a4[0]);
	assign C5j2a4 = (~(Hw63a4[0] | Hw63a4[1]));
	assign H4j2a4 = (~(Hw63a4[1] & J5j2a4));
	assign J5j2a4 = (Q5j2a4 | Hw63a4[0]);
	assign M3j2a4 = (Xx63a4[0] | Xx63a4[1]);
	assign F3j2a4 = (Hw63a4[0] | Hw63a4[1]);
	assign Lzi2a4 = (H1f2a4 & Bgb2a4);
	assign Bgb2a4 = (~(H1f2a4 & X5j2a4));
	assign H1f2a4 = (~(Js3x84 & E6j2a4));
	assign E6j2a4 = (~(L6j2a4 & X5j2a4));
	assign X5j2a4 = (S6j2a4 | V1f2a4);
	assign L6j2a4 = (~(Z6j2a4 & G7j2a4));
	assign G7j2a4 = (~(N7j2a4 & D373a4[0]));
	assign N7j2a4 = (~(K2j2a4 | U7j2a4));
	assign U7j2a4 = (D2j2a4 & B8j2a4);
	assign K2j2a4 = (V1f2a4 ? P8j2a4 : I8j2a4);
	assign Z6j2a4 = (B8j2a4 | D2j2a4);
	assign D2j2a4 = (V1f2a4 ? D9j2a4 : W8j2a4);
	assign V1f2a4 = (K9j2a4 & R9j2a4);
	assign R9j2a4 = (~(Y9j2a4 & S6j2a4));
	assign S6j2a4 = (~(G8i2a4 & Faj2a4));
	assign Faj2a4 = (~(K873a4[3] & R673a4[3]));
	assign Y9j2a4 = (~(Maj2a4 & Taj2a4));
	assign Taj2a4 = (~(Abj2a4 & D9j2a4));
	assign Maj2a4 = (Hbj2a4 | I8j2a4);
	assign I8j2a4 = (G8i2a4 ? Nz63a4[6] : Nz63a4[4]);
	assign Hbj2a4 = (~(P8j2a4 & Obj2a4));
	assign Obj2a4 = (D9j2a4 | Abj2a4);
	assign Abj2a4 = (!W8j2a4);
	assign P8j2a4 = (N8i2a4 ? Nz63a4[2] : Nz63a4[0]);
	assign K9j2a4 = (~(Vbj2a4 & N8i2a4));
	assign Vbj2a4 = (~(K873a4[1] & R673a4[1]));
	assign D9j2a4 = (N8i2a4 ? Nz63a4[3] : Nz63a4[1]);
	assign N8i2a4 = (~(Ccj2a4 & K873a4[0]));
	assign Ccj2a4 = (R673a4[0] & Jcj2a4);
	assign Jcj2a4 = (~(Qcj2a4 & Xcj2a4));
	assign Xcj2a4 = (Edj2a4 & Ldj2a4);
	assign Ldj2a4 = (~(Nz63a4[3] & Sdj2a4));
	assign Sdj2a4 = (~(Zdj2a4 & Nz63a4[0]));
	assign Zdj2a4 = (Nz63a4[1] & Gej2a4);
	assign Edj2a4 = (Nz63a4[1] | Nej2a4);
	assign Nej2a4 = (Nz63a4[0] & Gej2a4);
	assign Gej2a4 = (!Nz63a4[2]);
	assign Qcj2a4 = (K873a4[1] & R673a4[1]);
	assign W8j2a4 = (G8i2a4 ? Nz63a4[7] : Nz63a4[5]);
	assign G8i2a4 = (~(Uej2a4 & R673a4[2]));
	assign Uej2a4 = (K873a4[2] & Bfj2a4);
	assign Bfj2a4 = (~(Ifj2a4 & Pfj2a4));
	assign Pfj2a4 = (Wfj2a4 & Dgj2a4);
	assign Dgj2a4 = (~(Nz63a4[7] & Kgj2a4));
	assign Kgj2a4 = (Rgj2a4 | Ygj2a4);
	assign Wfj2a4 = (~(Ygj2a4 & Rgj2a4));
	assign Rgj2a4 = (!Nz63a4[5]);
	assign Ygj2a4 = (Fhj2a4 | Nz63a4[6]);
	assign Fhj2a4 = (!Nz63a4[4]);
	assign Ifj2a4 = (K873a4[3] & R673a4[3]);
	assign B8j2a4 = (!D373a4[1]);
	assign A1f2a4 = (~(Cc3x84 | La3x84));
	assign Cyi2a4 = (Mhj2a4 & Thj2a4);
	assign Thj2a4 = (~(Vlxx84 & V3ux84));
	assign Vlxx84 = (F5yx84 ? Q7yx84 : Kbyx84);
	assign Q7yx84 = (~(Aij2a4 & Hij2a4));
	assign Hij2a4 = (Oij2a4 & Vij2a4);
	assign Vij2a4 = (~(Htf2a4 & Sng2a4));
	assign Oij2a4 = (~(Aryx84 & Tkg2a4));
	assign Aij2a4 = (Cjj2a4 & Jjj2a4);
	assign Jjj2a4 = (~(Quf2a4 & Uog2a4));
	assign Cjj2a4 = (~(Tqyx84 & Vlg2a4));
	assign Kbyx84 = (~(Qjj2a4 & Xjj2a4));
	assign Xjj2a4 = (Ekj2a4 & Lkj2a4);
	assign Lkj2a4 = (~(Htf2a4 & Alg2a4));
	assign Ekj2a4 = (~(Aryx84 & Oeg2a4));
	assign Qjj2a4 = (Skj2a4 & Zkj2a4);
	assign Zkj2a4 = (~(Quf2a4 & Cmg2a4));
	assign Skj2a4 = (~(Tqyx84 & Qfg2a4));
	assign Mhj2a4 = (~(Pu63a4[15] & Pttx84));
	assign Oxi2a4 = (Glj2a4 & Nlj2a4);
	assign Nlj2a4 = (Ulj2a4 & Bmj2a4);
	assign Bmj2a4 = (~(X473a4[15] & Yutx84));
	assign Ulj2a4 = (~(HRDATA[15] & Fvtx84));
	assign Glj2a4 = (Imj2a4 & Pmj2a4);
	assign Pmj2a4 = (~(Nz63a4[3] & Awtx84));
	assign Imj2a4 = (~(STCALIB[15] & Hwtx84));
	assign Hxi2a4 = (Vx2x84 & Wmj2a4);
	assign Wmj2a4 = (Dnj2a4 | Vs63a4[1]);
	assign Twi2a4 = (~(Vs63a4[1] & Knj2a4));
	assign Knj2a4 = (~(Rnj2a4 & Ynj2a4));
	assign Ynj2a4 = (~(Foj2a4 & S9xx84));
	assign Foj2a4 = (~(Cmqx84 | Vs63a4[0]));
	assign Cmqx84 = (Moj2a4 & Toj2a4);
	assign Toj2a4 = (Apj2a4 & Hpj2a4);
	assign Hpj2a4 = (Opj2a4 & Vpj2a4);
	assign Vpj2a4 = (~(Pu63a4[23] & Pttx84));
	assign Pttx84 = (Cqj2a4 & R7hx84);
	assign Cqj2a4 = (Jqj2a4 & Scgx84);
	assign Opj2a4 = (~(X473a4[23] & Yutx84));
	assign Yutx84 = (Qqj2a4 & R7hx84);
	assign Qqj2a4 = (O3ux84 & Fhfx84);
	assign Fhfx84 = (Xqj2a4 & Q34x84);
	assign Xqj2a4 = (~(Wz3x84 | T14x84));
	assign Apj2a4 = (Erj2a4 & Lrj2a4);
	assign Lrj2a4 = (Snxx84 | Jve2a4);
	assign Jve2a4 = (!V3ux84);
	assign Snxx84 = (F5yx84 ? Xhe2a4 : H6yx84);
	assign Xhe2a4 = (Srj2a4 & Zrj2a4);
	assign Zrj2a4 = (Gsj2a4 & Nsj2a4);
	assign Nsj2a4 = (~(Htf2a4 & P4g2a4));
	assign Gsj2a4 = (~(Aryx84 & A7g2a4));
	assign Srj2a4 = (Usj2a4 & Btj2a4);
	assign Btj2a4 = (~(Quf2a4 & R5g2a4));
	assign Usj2a4 = (~(Tqyx84 & C8g2a4));
	assign H6yx84 = (Itj2a4 & Ptj2a4);
	assign Ptj2a4 = (Wtj2a4 & Duj2a4);
	assign Duj2a4 = (~(Htf2a4 & H7g2a4));
	assign Wtj2a4 = (~(Aryx84 & Lng2a4));
	assign Itj2a4 = (Kuj2a4 & Ruj2a4);
	assign Ruj2a4 = (~(Quf2a4 & J8g2a4));
	assign Kuj2a4 = (~(Tqyx84 & Nog2a4));
	assign Erj2a4 = (~(HRDATA[23] & Fvtx84));
	assign Moj2a4 = (Yuj2a4 & Fvj2a4);
	assign Fvj2a4 = (~(STCALIB[23] & Hwtx84));
	assign Yuj2a4 = (Mvj2a4 & Tvj2a4);
	assign Tvj2a4 = (~(W0ux84 & Hw63a4[1]));
	assign Mvj2a4 = (~(Nz63a4[5] & Awtx84));
	assign Rnj2a4 = (Dnj2a4 | Hlqx84);
	assign Hlqx84 = (Awj2a4 & Hwj2a4);
	assign Hwj2a4 = (Owj2a4 & Vwj2a4);
	assign Vwj2a4 = (Cxj2a4 & Jxj2a4);
	assign Jxj2a4 = (~(Qxj2a4 & Cahx84));
	assign Cahx84 = (Xxj2a4 & Eyj2a4);
	assign Xxj2a4 = (V2hx84 & T14x84);
	assign Qxj2a4 = (Xx63a4[1] & O3ux84);
	assign Cxj2a4 = (Hge2a4 & Lyj2a4);
	assign Lyj2a4 = (!Vge2a4);
	assign Vge2a4 = (Woyx84 & V3ux84);
	assign Woyx84 = (!Luxx84);
	assign Luxx84 = (~(Syj2a4 & Zyj2a4));
	assign Zyj2a4 = (Gzj2a4 & F7bx84);
	assign Gzj2a4 = (Atix84 & K5g2a4);
	assign Syj2a4 = (Me5w84 & Ub82a4);
	assign Hge2a4 = (~(Nzj2a4 & Uzj2a4));
	assign Uzj2a4 = (Eyj2a4 & I6hx84);
	assign Eyj2a4 = (~(Scgx84 | Wz3x84));
	assign Nzj2a4 = (T14x84 & O3ux84);
	assign Owj2a4 = (B0k2a4 & I0k2a4);
	assign I0k2a4 = (~(La3x84 & Gstx84));
	assign Gstx84 = (O3ux84 & Wpjx84);
	assign Wpjx84 = (Z9g2a4 & I6hx84);
	assign Z9g2a4 = (P0k2a4 & Q34x84);
	assign P0k2a4 = (~(Dfgx84 | T14x84));
	assign B0k2a4 = (~(Uvxx84 & V3ux84));
	assign V3ux84 = (Me5w84 & W0k2a4);
	assign W0k2a4 = (~(D1k2a4 & K1k2a4));
	assign K1k2a4 = (~(O8px84 | Yzhx84));
	assign D1k2a4 = (R1k2a4 & Y1k2a4);
	assign Y1k2a4 = (Mmvx84 | J13x84);
	assign R1k2a4 = (Qxmx84 | Ns2x84);
	assign Uvxx84 = (~(Iye2a4 | Xmxx84));
	assign Xmxx84 = (F5yx84 ? Vkyx84 : Eie2a4);
	assign Vkyx84 = (F2k2a4 & M2k2a4);
	assign M2k2a4 = (T2k2a4 & A3k2a4);
	assign A3k2a4 = (~(Htf2a4 & Ixf2a4));
	assign T2k2a4 = (~(Aryx84 & Otf2a4));
	assign F2k2a4 = (H3k2a4 & O3k2a4);
	assign O3k2a4 = (~(Quf2a4 & Kyf2a4));
	assign H3k2a4 = (~(Tqyx84 & Xuf2a4));
	assign Eie2a4 = (V3k2a4 & C4k2a4);
	assign C4k2a4 = (J4k2a4 & Q4k2a4);
	assign Q4k2a4 = (~(Htf2a4 & Vtf2a4));
	assign Htf2a4 = (~(X4k2a4 | E5k2a4));
	assign J4k2a4 = (~(Aryx84 & I4g2a4));
	assign Aryx84 = (X4k2a4 & L5k2a4);
	assign V3k2a4 = (S5k2a4 & Z5k2a4);
	assign Z5k2a4 = (~(Quf2a4 & Evf2a4));
	assign Quf2a4 = (G6k2a4 & E5k2a4);
	assign G6k2a4 = (!X4k2a4);
	assign S5k2a4 = (~(Tqyx84 & K5g2a4));
	assign Iye2a4 = (~(Hryx84 & N6k2a4));
	assign N6k2a4 = (Pye2a4 | F5h2a4);
	assign F5h2a4 = (!Tqyx84);
	assign Pye2a4 = (!Fqyx84);
	assign Fqyx84 = (U6k2a4 & Wbcx84);
	assign U6k2a4 = (~(Aff2a4 ^ F5yx84));
	assign Hryx84 = (~(B7k2a4 & Aff2a4));
	assign Aff2a4 = (!K4h2a4);
	assign K4h2a4 = (~(Zfyx84 | I7k2a4));
	assign Zfyx84 = (!Ugyx84);
	assign Ugyx84 = (~(Rybx84 & P7k2a4));
	assign P7k2a4 = (Zo2x84 | Bw2x84);
	assign B7k2a4 = (~(Tqyx84 | Wlnx84));
	assign Awj2a4 = (W7k2a4 & D8k2a4);
	assign D8k2a4 = (K8k2a4 & R8k2a4);
	assign R8k2a4 = (~(HRDATA[31] & Fvtx84));
	assign Fvtx84 = (S9g2a4 & J0kx84);
	assign J0kx84 = (Y8k2a4 & Dfgx84);
	assign Dfgx84 = (!Wz3x84);
	assign S9g2a4 = (V2hx84 & O3ux84);
	assign V2hx84 = (~(Cw3x84 | Zx3x84));
	assign K8k2a4 = (~(W0ux84 & D373a4[1]));
	assign W0ux84 = (F9k2a4 & Jqj2a4);
	assign F9k2a4 = (I6hx84 & Scgx84);
	assign Scgx84 = (!Q34x84);
	assign I6hx84 = (Zx3x84 & Vjex84);
	assign W7k2a4 = (M9k2a4 & T9k2a4);
	assign T9k2a4 = (~(Nz63a4[7] & Awtx84));
	assign Awtx84 = (Aak2a4 & M8hx84);
	assign M8hx84 = (Y8k2a4 & Wz3x84);
	assign Y8k2a4 = (~(T14x84 | Q34x84));
	assign Aak2a4 = (O3ux84 & T8hx84);
	assign T8hx84 = (Cw3x84 & Zx3x84);
	assign M9k2a4 = (~(STCALIB[25] & Hwtx84));
	assign Hwtx84 = (Hak2a4 & R7hx84);
	assign R7hx84 = (~(Vjex84 | Zx3x84));
	assign Vjex84 = (!Cw3x84);
	assign Hak2a4 = (Jqj2a4 & Q34x84);
	assign Jqj2a4 = (Oak2a4 & T14x84);
	assign Oak2a4 = (O3ux84 & Wz3x84);
	assign Dnj2a4 = (Hu2x84 & Vak2a4);
	assign Vak2a4 = (~(Vs63a4[0] & S9xx84));
	assign S9xx84 = (Mgnx84 & G4bx84);
	assign Hhux84 = (Rprx84 & Lfyx84);
	assign Lfyx84 = (M0wx84 | Ufi2a4);
	assign Ufi2a4 = (Wpxx84 & Cbk2a4);
	assign Cbk2a4 = (!I7k2a4);
	assign I7k2a4 = (Jbk2a4 & Tqyx84);
	assign Tqyx84 = (E5k2a4 & X4k2a4);
	assign X4k2a4 = (Qbk2a4 | Xbk2a4);
	assign Qbk2a4 = (Lck2a4 ? Eck2a4 : Fkxx84);
	assign Eck2a4 = (~(E5k2a4 | Fkxx84));
	assign Jbk2a4 = (~(Sck2a4 | F5yx84));
	assign F5yx84 = (!Gxe2a4);
	assign Gxe2a4 = (~(Zck2a4 & Gdk2a4));
	assign Zck2a4 = (Wpxx84 ? Udk2a4 : Ndk2a4);
	assign Udk2a4 = (~(Bek2a4 & Ndk2a4));
	assign Sck2a4 = (!Yqxx84);
	assign M0wx84 = (!Nvxx84);
	assign Nvxx84 = (Yqxx84 & Xlyx84);
	assign Xlyx84 = (Wlnx84 | Iixx84);
	assign Iixx84 = (Iek2a4 & Pek2a4);
	assign Pek2a4 = (Wek2a4 | Dfk2a4);
	assign Iek2a4 = (Bpxx84 & Kfk2a4);
	assign Kfk2a4 = (~(Rfk2a4 & Yfk2a4));
	assign Yfk2a4 = (Fgk2a4 & Itmx84);
	assign Fgk2a4 = (~(Ap6w84 | Zo2x84));
	assign Rfk2a4 = (Mgk2a4 & Tgk2a4);
	assign Mgk2a4 = (~(Evix84 | Wl6w84));
	assign Bpxx84 = (~(Ahk2a4 & Hhk2a4));
	assign Hhk2a4 = (~(Ohk2a4 & Vhk2a4));
	assign Yqxx84 = (~(Osxx84 | Olxx84));
	assign Olxx84 = (Cik2a4 & Ipxx84);
	assign Ipxx84 = (Jik2a4 | Qik2a4);
	assign Cik2a4 = (Fkxx84 ? Qik2a4 : Xik2a4);
	assign Fkxx84 = (!Wpxx84);
	assign Xik2a4 = (~(Qik2a4 & Jik2a4));
	assign Qik2a4 = (~(Ejk2a4 & Ljk2a4));
	assign Ljk2a4 = (Sjk2a4 | Wek2a4);
	assign Ejk2a4 = (D8gx84 | Evix84);
	assign Osxx84 = (!Cmxx84);
	assign Cmxx84 = (~(Zjk2a4 & Jik2a4));
	assign Jik2a4 = (Gdk2a4 | Gkk2a4);
	assign Zjk2a4 = (Wpxx84 ? Nkk2a4 : Gkk2a4);
	assign Wpxx84 = (~(Rybx84 & Ukk2a4));
	assign Ukk2a4 = (O8bx84 | Bw2x84);
	assign Nkk2a4 = (~(Gkk2a4 & Gdk2a4));
	assign Gdk2a4 = (Ndk2a4 | Bek2a4);
	assign Bek2a4 = (!Xbk2a4);
	assign Xbk2a4 = (Blk2a4 & E5k2a4);
	assign E5k2a4 = (!L5k2a4);
	assign L5k2a4 = (~(Ilk2a4 & Plk2a4));
	assign Plk2a4 = (Wlk2a4 | Wek2a4);
	assign Ilk2a4 = (Tn1y84 | Evix84);
	assign Blk2a4 = (!Lck2a4);
	assign Lck2a4 = (~(Dmk2a4 & Kmk2a4));
	assign Kmk2a4 = (Rmk2a4 | Wek2a4);
	assign Dmk2a4 = (Hanx84 | Evix84);
	assign Ndk2a4 = (~(Ymk2a4 & Fnk2a4));
	assign Fnk2a4 = (Mnk2a4 | Wek2a4);
	assign Wek2a4 = (!Ahk2a4);
	assign Ymk2a4 = (Bf0y84 | Evix84);
	assign Gkk2a4 = (~(Tnk2a4 & Aok2a4));
	assign Aok2a4 = (~(Hok2a4 & Ahk2a4));
	assign Ahk2a4 = (~(K2c2a4 & Ny1y84));
	assign Ny1y84 = (!C0dx84);
	assign C0dx84 = (Hu2x84 & Tsix84);
	assign K2c2a4 = (O8bx84 | Ewax84);
	assign Tnk2a4 = (Itmx84 | Evix84);
	assign Gmi2a4 = (Pvrx84 | Rprx84);
	assign Rprx84 = (!Orrx84);
	assign Orrx84 = (~(Ook2a4 & Vok2a4));
	assign Vok2a4 = (~(Cpk2a4 & Axb2a4));
	assign Cpk2a4 = (J13x84 | Mlbx84);
	assign Ook2a4 = (Jpk2a4 & Dybx84);
	assign Jpk2a4 = (~(Atix84 & Qpk2a4));
	assign Qpk2a4 = (Qxmx84 | Drbx84);
	assign Pvrx84 = (~(HRESP & O3ux84));
	assign O3ux84 = (Me5w84 & Xpk2a4);
	assign Xpk2a4 = (~(Eqk2a4 & Lqk2a4));
	assign Lqk2a4 = (Sqk2a4 & Ambx84);
	assign Sqk2a4 = (~(Zqk2a4 & Zvix84));
	assign Zqk2a4 = (~(Ewax84 | Hu2x84));
	assign Eqk2a4 = (Grk2a4 & Nrk2a4);
	assign Nrk2a4 = (~(Urk2a4 & Uacx84));
	assign Urk2a4 = (~(Xtcx84 | Fn2x84));
	assign Xtcx84 = (!Atix84);
	assign Grk2a4 = (~(Mlbx84 & H6dx84));
	assign F8e2a4 = (~(T0wx84 & Nocx84));
	assign T0wx84 = (Mrcx84 & Gcvx84);
	assign Mrcx84 = (Tq2x84 & G4bx84);
	assign Xlh2a4 = (~(Qoe2a4 & Es0x84));
	assign Qoe2a4 = (Acex84 & Dj0x84);
	assign Acex84 = (Nocx84 & Bsk2a4);
	assign Bsk2a4 = (~(Fbex84 & Isk2a4));
	assign Isk2a4 = (F2gx84 | Mbex84);
	assign Fbex84 = (Tq2x84 & Ewax84);
	assign Nocx84 = (HREADY & Hscx84);
	assign Hscx84 = (~(Psk2a4 & Wsk2a4));
	assign Wsk2a4 = (Dtk2a4 & Ktk2a4);
	assign Ktk2a4 = (~(Rtk2a4 & N4ix84));
	assign Rtk2a4 = (~(Yqcx84 | T7bx84));
	assign Dtk2a4 = (~(Wlnx84 & Ytk2a4));
	assign Ytk2a4 = (~(Fuk2a4 & Muk2a4));
	assign Muk2a4 = (Jxmx84 | Tswx84);
	assign Fuk2a4 = (~(Nwix84 & Uj2x84));
	assign Psk2a4 = (Ylvx84 & Tuk2a4);
	assign Tuk2a4 = (F5dx84 | Lrfx84);
	assign Ylvx84 = (Gqox84 | Fn2x84);
	assign Xaax84 = (~(Avk2a4 ^ Slzx84));
	assign Avk2a4 = (~(Hvk2a4 & Ovk2a4));
	assign Ovk2a4 = (Sr0y84 | Kozx84);
	assign Hvk2a4 = (Vvk2a4 & Tpzx84);
	assign Vvk2a4 = (~(Tt6w84 & Dozx84));
	assign Qaax84 = (~(Cwk2a4 ^ Slzx84));
	assign Cwk2a4 = (~(Jwk2a4 & Qwk2a4));
	assign Qwk2a4 = (Du0y84 | Kozx84);
	assign Jwk2a4 = (Xwk2a4 & Tpzx84);
	assign Xwk2a4 = (~(Iv6w84 & Dozx84));
	assign Jaax84 = (~(Exk2a4 ^ Slzx84));
	assign Exk2a4 = (~(Lxk2a4 & Sxk2a4));
	assign Sxk2a4 = (B01y84 | Kozx84);
	assign Lxk2a4 = (Zxk2a4 & Tpzx84);
	assign Zxk2a4 = (~(Hk6w84 & Dozx84));
	assign Caax84 = (~(Gyk2a4 ^ Slzx84));
	assign Gyk2a4 = (~(Nyk2a4 & Uyk2a4));
	assign Uyk2a4 = (Nd1y84 | Kozx84);
	assign Nyk2a4 = (Bzk2a4 & Tpzx84);
	assign Bzk2a4 = (~(Es6w84 & Dozx84));
	assign V9ax84 = (W8tx84 ? Axzx84 : Hxzx84);
	assign O9ax84 = (Yf1y84 ? Hxzx84 : Axzx84);
	assign H9ax84 = (Dwdx84 ? Axzx84 : Hxzx84);
	assign A9ax84 = (Vitx84 ? Axzx84 : Hxzx84);
	assign Axzx84 = (X50y84 | E60y84);
	assign E60y84 = (Slzx84 & Izk2a4);
	assign X50y84 = (Pzk2a4 | Wzk2a4);
	assign Wzk2a4 = (Kozx84 & L60y84);
	assign Hxzx84 = (Pzk2a4 | L60y84);
	assign L60y84 = (D0l2a4 & Tpzx84);
	assign D0l2a4 = (~(W10y84 | Slzx84));
	assign Pzk2a4 = (Slzx84 & K0l2a4);
	assign K0l2a4 = (~(Tpzx84 & Qyzx84));
	assign Qyzx84 = (!W10y84);
	assign W10y84 = (C07w84 & Dozx84);
	assign Tpzx84 = (Fwzx84 | T7px84);
	assign T8ax84 = (~(R0l2a4 ^ Slzx84));
	assign R0l2a4 = (~(Y0l2a4 & F1l2a4));
	assign F1l2a4 = (M1l2a4 & T1l2a4);
	assign T1l2a4 = (~(Es6w84 & Inzx84));
	assign M1l2a4 = (~(G36w84 & Dozx84));
	assign Y0l2a4 = (A2l2a4 & H2l2a4);
	assign H2l2a4 = (Dnmx84 | Fwzx84);
	assign A2l2a4 = (M21y84 | Kozx84);
	assign M8ax84 = (~(O2l2a4 ^ Slzx84));
	assign O2l2a4 = (~(V2l2a4 & C3l2a4));
	assign C3l2a4 = (J3l2a4 & Q3l2a4);
	assign Q3l2a4 = (~(Es6w84 & Bnzx84));
	assign J3l2a4 = (~(Inzx84 & Ap6w84));
	assign V2l2a4 = (X3l2a4 & E4l2a4);
	assign E4l2a4 = (~(Dozx84 & Wz5w84));
	assign X3l2a4 = (X41y84 | Kozx84);
	assign F8ax84 = (~(L4l2a4 ^ Slzx84));
	assign L4l2a4 = (~(S4l2a4 & Z4l2a4));
	assign Z4l2a4 = (G5l2a4 & N5l2a4);
	assign N5l2a4 = (Itmx84 | Gl0y84);
	assign Itmx84 = (!Ln6w84);
	assign G5l2a4 = (~(Pq6w84 & Bnzx84));
	assign S4l2a4 = (U5l2a4 & B6l2a4);
	assign B6l2a4 = (~(Dozx84 & Ey5w84));
	assign U5l2a4 = (Vw0y84 | Kozx84);
	assign Y7ax84 = (~(I6l2a4 ^ Slzx84));
	assign I6l2a4 = (~(P6l2a4 & W6l2a4));
	assign W6l2a4 = (D7l2a4 & K7l2a4);
	assign K7l2a4 = (Bf0y84 | Gl0y84);
	assign Gl0y84 = (~(Inzx84 | R7l2a4));
	assign R7l2a4 = (Ol2x84 & Y7l2a4);
	assign Y7l2a4 = (~(F8l2a4 & M8l2a4));
	assign M8l2a4 = (~(T8l2a4 | L3ix84));
	assign L3ix84 = (J13x84 & Ns2x84);
	assign T8l2a4 = (Dzox84 | Iqbx84);
	assign Dzox84 = (E3wx84 & Y6bx84);
	assign F8l2a4 = (Cldx84 & A9l2a4);
	assign A9l2a4 = (Cuix84 | Vx2x84);
	assign Cuix84 = (!E3wx84);
	assign Cldx84 = (~(Aq42a4 | Frcx84));
	assign Bf0y84 = (!Wl6w84);
	assign D7l2a4 = (~(Ap6w84 & Bnzx84));
	assign Bnzx84 = (~(H9l2a4 & O9l2a4));
	assign O9l2a4 = (~(I5bx84 & V9l2a4));
	assign V9l2a4 = (~(Cal2a4 & Jal2a4));
	assign Jal2a4 = (Tsix84 | Vx2x84);
	assign Cal2a4 = (Qal2a4 & Xal2a4);
	assign Xal2a4 = (M6xx84 | Bs1y84);
	assign M6xx84 = (!Gpix84);
	assign Qal2a4 = (Bdox84 | F5dx84);
	assign H9l2a4 = (Ebl2a4 & Fwzx84);
	assign Ebl2a4 = (~(Ol2x84 & Lbl2a4));
	assign Lbl2a4 = (~(Sbl2a4 & Zbl2a4));
	assign Zbl2a4 = (~(Gcl2a4 & J982a4));
	assign Gcl2a4 = (Pz2x84 & U4px84);
	assign U4px84 = (Yqcx84 | Gz4w84);
	assign Sbl2a4 = (~(Ncl2a4 & Tq2x84));
	assign Ncl2a4 = (Ucl2a4 & Ambx84);
	assign Ucl2a4 = (~(Kshx84 & Bdl2a4));
	assign Bdl2a4 = (S1dx84 | Vx2x84);
	assign Kshx84 = (!Y6bx84);
	assign P6l2a4 = (Idl2a4 & Pdl2a4);
	assign Pdl2a4 = (~(Mw5w84 & Dozx84));
	assign Idl2a4 = (W71y84 | Kozx84);
	assign R7ax84 = (~(Wdl2a4 ^ Slzx84));
	assign Slzx84 = (Del2a4 & Kel2a4);
	assign Kel2a4 = (~(I5bx84 & Rel2a4));
	assign Rel2a4 = (~(Yel2a4 & Ffl2a4));
	assign Ffl2a4 = (~(Mfl2a4 & Yzhx84));
	assign Mfl2a4 = (~(O8bx84 | Ewax84));
	assign Yel2a4 = (Mycx84 | Tsix84);
	assign Del2a4 = (Xvax84 | Tfl2a4);
	assign Tfl2a4 = (Agl2a4 & V8bx84);
	assign V8bx84 = (Hgl2a4 & Ogl2a4);
	assign Ogl2a4 = (Fycx84 | Evix84);
	assign Hgl2a4 = (Vgl2a4 & Chl2a4);
	assign Chl2a4 = (~(Jhl2a4 & E3wx84));
	assign Jhl2a4 = (Laix84 & Y3i2a4);
	assign Vgl2a4 = (Bs1y84 | F5dx84);
	assign Bs1y84 = (!Klvx84);
	assign Agl2a4 = (Qhl2a4 & Xhl2a4);
	assign Xhl2a4 = (~(Pz2x84 & Eil2a4));
	assign Eil2a4 = (~(Lil2a4 & Sil2a4));
	assign Sil2a4 = (Sbox84 | Gpbx84);
	assign Sbox84 = (!Mbex84);
	assign Mbex84 = (Zo2x84 & G4bx84);
	assign Lil2a4 = (Qw1y84 | Fycx84);
	assign Wdl2a4 = (~(Zil2a4 & Gjl2a4));
	assign Gjl2a4 = (Njl2a4 & Ujl2a4);
	assign Ujl2a4 = (~(Inzx84 & Tt6w84));
	assign Inzx84 = (Ol2x84 & Bkl2a4);
	assign Bkl2a4 = (~(Ikl2a4 & Pkl2a4));
	assign Pkl2a4 = (Wkl2a4 & T7bx84);
	assign T7bx84 = (V2ox84 | Mmvx84);
	assign Wkl2a4 = (~(Dll2a4 & Sz42a4));
	assign Dll2a4 = (~(Qw1y84 | J13x84));
	assign Ikl2a4 = (Kll2a4 & Rll2a4);
	assign Rll2a4 = (~(Gz4w84 & Yll2a4));
	assign Yll2a4 = (~(Uy1y84 & Fml2a4));
	assign Fml2a4 = (~(Mml2a4 & G4bx84));
	assign Mml2a4 = (Lw72a4 | Y6bx84);
	assign Kll2a4 = (Mzbx84 | Wqbx84);
	assign Mzbx84 = (!Teix84);
	assign Teix84 = (J13x84 & Yqcx84);
	assign Njl2a4 = (~(Y46w84 & Dozx84));
	assign Dozx84 = (Tml2a4 & Jm92a4);
	assign Tml2a4 = (~(Ebox84 | Xvax84));
	assign Ebox84 = (!O1px84);
	assign O1px84 = (Hu2x84 & Yqcx84);
	assign Zil2a4 = (Anl2a4 & Hnl2a4);
	assign Hnl2a4 = (Kkbx84 | Fwzx84);
	assign Fwzx84 = (~(Onl2a4 & Vnl2a4));
	assign Onl2a4 = (~(Xvax84 | H8px84));
	assign Kkbx84 = (!Xw6w84);
	assign Anl2a4 = (Cb1y84 | Kozx84);
	assign Kozx84 = (!Izk2a4);
	assign Izk2a4 = (~(Col2a4 & Jol2a4));
	assign Jol2a4 = (~(I5bx84 & Qol2a4));
	assign Qol2a4 = (~(W1c2a4 & Xol2a4));
	assign Xol2a4 = (Fmvx84 | Bw2x84);
	assign I5bx84 = (~(Xvax84 | Pz2x84));
	assign Xvax84 = (!Ol2x84);
	assign Col2a4 = (~(Ol2x84 & Epl2a4));
	assign Epl2a4 = (~(Lpl2a4 & Spl2a4));
	assign Spl2a4 = (~(Ja72a4 | Nndx84));
	assign Ja72a4 = (Zpl2a4 & Gcvx84);
	assign Zpl2a4 = (~(Qxmx84 | Ns2x84));
	assign Lpl2a4 = (Gql2a4 & Nql2a4);
	assign Nql2a4 = (~(Uql2a4 & F2gx84));
	assign Uql2a4 = (~(Dybx84 | Hu2x84));
	assign Gql2a4 = (~(Gz4w84 & Brl2a4));
	assign Brl2a4 = (~(Irl2a4 & Prl2a4));
	assign Prl2a4 = (~(Dt62a4 & Fn2x84));
	assign Dt62a4 = (~(Tq2x84 | Bw2x84));
	assign Irl2a4 = (O8bx84 | Ns2x84);
	assign O8bx84 = (!Uwix84);
	assign TXEV = (Wrl2a4 & Y6bx84);
	assign Wrl2a4 = (~(Gpbx84 | Mmvx84));
	assign SLEEPDEEP = (SLEEPING & Y63x84);
	assign SLEEPING = (Bh3x84 & Tbex84);
	assign Tbex84 = (!Ju4w84);
	assign LOCKUP = (~(Dsl2a4 & Ksl2a4));
	assign Ksl2a4 = (Rsl2a4 | Ambx84);
	assign Dsl2a4 = (Ysl2a4 & Ftl2a4);
	assign Ftl2a4 = (~(Mtl2a4 & Sz42a4));
	assign Sz42a4 = (~(H8px84 | D4dx84));
	assign Mtl2a4 = (Vnl2a4 & Qxmx84);
	assign Ysl2a4 = (~(G33x84 & Ttl2a4));
	assign Ttl2a4 = (~(Mblx84 & Aul2a4));
	assign Aul2a4 = (~(Oclx84 & Ns2x84));
	assign Oclx84 = (Hul2a4 & Hx42a4);
	assign Hul2a4 = (Tamx84 & Rv42a4);
	assign Mblx84 = (Oul2a4 & Vul2a4);
	assign Vul2a4 = (Cvl2a4 & Jvl2a4);
	assign Jvl2a4 = (~(Lb2y84 & Qvl2a4));
	assign Qvl2a4 = (Tamx84 & Vx2x84);
	assign Lb2y84 = (~(A0cx84 | N4bx84));
	assign Cvl2a4 = (Xvl2a4 & Ewl2a4);
	assign Xvl2a4 = (~(Lwl2a4 & Swl2a4));
	assign Swl2a4 = (Zwl2a4 & Hgvx84);
	assign Zwl2a4 = (~(Gxl2a4 & Yv42a4));
	assign Yv42a4 = (!Hx42a4);
	assign Hx42a4 = (B9lx84 & Gpix84);
	assign Gxl2a4 = (~(Auox84 & Ykwx84));
	assign Ykwx84 = (Ub82a4 & Jm92a4);
	assign Auox84 = (~(Ns2x84 | Hu2x84));
	assign Lwl2a4 = (~(T692a4 | Nxl2a4));
	assign Nxl2a4 = (~(F3mx84 | Jtcx84));
	assign Oul2a4 = (Uxl2a4 & Byl2a4);
	assign Byl2a4 = (Iyl2a4 | B5bx84);
	assign Uxl2a4 = (Pyl2a4 & Wyl2a4);
	assign Wyl2a4 = (~(Dzl2a4 & Kikx84));
	assign Kikx84 = (~(A0cx84 | P1mx84));
	assign A0cx84 = (!Jm92a4);
	assign Dzl2a4 = (~(Qxmx84 | Ssex84));
	assign Ssex84 = (!Phkx84);
	assign Phkx84 = (~(Kzl2a4 & Rzl2a4));
	assign Rzl2a4 = (~(Yzl2a4 & P8c2a4));
	assign P8c2a4 = (~(F0m2a4 & M0m2a4));
	assign M0m2a4 = (T0m2a4 & A1m2a4);
	assign A1m2a4 = (~(Nojx84 | Ihkx84));
	assign T0m2a4 = (~(Yqjx84 | Dlhx84));
	assign F0m2a4 = (H1m2a4 & Y9fx84);
	assign Y9fx84 = (!X0kx84);
	assign H1m2a4 = (~(Umex84 | Ctjx84));
	assign Yzl2a4 = (~(O1m2a4 & V1m2a4));
	assign V1m2a4 = (~(Xx63a4[1] & C2m2a4));
	assign C2m2a4 = (J2m2a4 | G7c2a4);
	assign O1m2a4 = (~(G7c2a4 & J2m2a4));
	assign J2m2a4 = (~(Q5j2a4 & Z6c2a4));
	assign Z6c2a4 = (~(Q2m2a4 & X2m2a4));
	assign X2m2a4 = (E3m2a4 & L3m2a4);
	assign L3m2a4 = (S3m2a4 & Z3m2a4);
	assign Z3m2a4 = (~(Nz63a4[4] & Yqjx84));
	assign S3m2a4 = (~(Nz63a4[6] & X0kx84));
	assign E3m2a4 = (G4m2a4 & N4m2a4);
	assign N4m2a4 = (~(Nz63a4[2] & Ctjx84));
	assign G4m2a4 = (~(Nz63a4[0] & Umex84));
	assign Q2m2a4 = (U4m2a4 & B5m2a4);
	assign B5m2a4 = (~(Ihkx84 & Xx63a4[0]));
	assign U4m2a4 = (I5m2a4 & P5m2a4);
	assign P5m2a4 = (~(Dlhx84 & Hw63a4[0]));
	assign I5m2a4 = (~(Nojx84 & D373a4[0]));
	assign Q5j2a4 = (!Xx63a4[0]);
	assign G7c2a4 = (W5m2a4 & D6m2a4);
	assign D6m2a4 = (K6m2a4 & R6m2a4);
	assign R6m2a4 = (Y6m2a4 & F7m2a4);
	assign F7m2a4 = (~(Nz63a4[5] & Yqjx84));
	assign Yqjx84 = (M7m2a4 & T7m2a4);
	assign M7m2a4 = (~(Omf2a4 | Nj63a4[0]));
	assign Y6m2a4 = (~(Nz63a4[7] & X0kx84));
	assign X0kx84 = (A8m2a4 & Nj63a4[0]);
	assign A8m2a4 = (T7m2a4 & Nj63a4[1]);
	assign K6m2a4 = (H8m2a4 & O8m2a4);
	assign O8m2a4 = (~(Nz63a4[3] & Ctjx84));
	assign Ctjx84 = (V8m2a4 & Nj63a4[0]);
	assign V8m2a4 = (T7m2a4 & Omf2a4);
	assign H8m2a4 = (~(Nz63a4[1] & Umex84));
	assign Umex84 = (C9m2a4 & T7m2a4);
	assign T7m2a4 = (J9m2a4 & Q9m2a4);
	assign Q9m2a4 = (~(Nj63a4[3] | Nj63a4[5]));
	assign J9m2a4 = (Nj63a4[4] & Rqg2a4);
	assign C9m2a4 = (~(Nj63a4[0] | Nj63a4[1]));
	assign W5m2a4 = (X9m2a4 & Eam2a4);
	assign Eam2a4 = (~(Ihkx84 & Xx63a4[1]));
	assign Ihkx84 = (Lam2a4 & Sam2a4);
	assign Lam2a4 = (~(Tbb2a4 | Nj63a4[2]));
	assign X9m2a4 = (Zam2a4 & Gbm2a4);
	assign Gbm2a4 = (~(Dlhx84 & Hw63a4[1]));
	assign Dlhx84 = (Nbm2a4 & Sam2a4);
	assign Nbm2a4 = (~(Rqg2a4 | Nj63a4[0]));
	assign Zam2a4 = (~(Nojx84 & D373a4[1]));
	assign Nojx84 = (Ubm2a4 & Sam2a4);
	assign Sam2a4 = (Bcm2a4 & Icm2a4);
	assign Bcm2a4 = (~(K7e2a4 | Omf2a4));
	assign Ubm2a4 = (~(Rqg2a4 | Tbb2a4));
	assign Rqg2a4 = (!Nj63a4[2]);
	assign Kzl2a4 = (~(Dmux84 | Nr4w84));
	assign Dmux84 = (!E7lx84);
	assign E7lx84 = (~(Pcm2a4 & Wcm2a4));
	assign Pcm2a4 = (~(Omf2a4 | Nj63a4[2]));
	assign Omf2a4 = (!Nj63a4[1]);
	assign Pyl2a4 = (~(Ddm2a4 & D53x84));
	assign Ddm2a4 = (~(Gpbx84 | Zo2x84));
	assign HWRITE = (~(Kdm2a4 & Rdm2a4));
	assign Rdm2a4 = (Ydm2a4 & Gqox84);
	assign Ydm2a4 = (Qnix84 & Fem2a4);
	assign Qnix84 = (~(Qvax84 & Lw72a4));
	assign Kdm2a4 = (Mem2a4 & Tem2a4);
	assign Tem2a4 = (~(Afm2a4 & Mmvx84));
	assign Afm2a4 = (~(Hfm2a4 & Ofm2a4));
	assign Ofm2a4 = (~(Vfm2a4 & Frcx84));
	assign Frcx84 = (Gcvx84 & Xm92a4);
	assign Vfm2a4 = (~(Qw1y84 | N4ix84));
	assign Qw1y84 = (!O8px84);
	assign O8px84 = (Fn2x84 & Hu2x84);
	assign Hfm2a4 = (Y4dx84 | Bdox84);
	assign Y4dx84 = (!Gc72a4);
	assign Mem2a4 = (Cgm2a4 & Jgm2a4);
	assign Jgm2a4 = (~(Qgm2a4 & Wyox84));
	assign Wyox84 = (J982a4 & Wqbx84);
	assign Qgm2a4 = (~(N4ix84 | Vx2x84));
	assign Cgm2a4 = (~(Xgm2a4 & Gc72a4));
	assign Xgm2a4 = (~(N4bx84 | Jnix84));
	assign HWDATA[9] = (!M3fx84);
	assign M3fx84 = (Ehm2a4 ? Sd0y84 : Cb1y84);
	assign HWDATA[8] = (!Lhm2a4);
	assign Lhm2a4 = (Ehm2a4 ? Yn0y84 : M21y84);
	assign HWDATA[7] = (C45w84 & Mizx84);
	assign HWDATA[6] = (~(Ralx84 | X41y84));
	assign HWDATA[5] = (~(Ralx84 | Vw0y84));
	assign HWDATA[4] = (C45w84 & Shm2a4);
	assign HWDATA[3] = (~(Ralx84 | Tlpx84));
	assign HWDATA[31] = (~(Zhm2a4 & Gim2a4));
	assign Gim2a4 = (Nim2a4 | Piqx84);
	assign Zhm2a4 = (Uim2a4 & Bjm2a4);
	assign Bjm2a4 = (~(N8b2a4 & Ysvx84));
	assign Ysvx84 = (~(Ijm2a4 & Pjm2a4));
	assign Pjm2a4 = (Wjm2a4 & Dkm2a4);
	assign Dkm2a4 = (Kkm2a4 & Rkm2a4);
	assign Rkm2a4 = (Ykm2a4 & Flm2a4);
	assign Flm2a4 = (~(S0hw84 & Mlm2a4));
	assign Ykm2a4 = (Tlm2a4 & Amm2a4);
	assign Amm2a4 = (~(Kwyw84 & Hmm2a4));
	assign Tlm2a4 = (~(Mf0x84 & Omm2a4));
	assign Kkm2a4 = (Vmm2a4 & Cnm2a4);
	assign Cnm2a4 = (~(Yhaw84 & Jnm2a4));
	assign Vmm2a4 = (~(Kniw84 & Qnm2a4));
	assign Wjm2a4 = (Xnm2a4 & Eom2a4);
	assign Eom2a4 = (Lom2a4 & Som2a4);
	assign Som2a4 = (~(Q4cw84 & Zom2a4));
	assign Lom2a4 = (~(Irdw84 & Gpm2a4));
	assign Xnm2a4 = (Npm2a4 & Upm2a4);
	assign Upm2a4 = (~(Cakw84 & Bqm2a4));
	assign Npm2a4 = (~(Aefw84 & Iqm2a4));
	assign Ijm2a4 = (Pqm2a4 & Wqm2a4);
	assign Wqm2a4 = (Drm2a4 & Krm2a4);
	assign Krm2a4 = (Rrm2a4 & Yrm2a4);
	assign Yrm2a4 = (~(Uwlw84 & Fsm2a4));
	assign Rrm2a4 = (~(Mjnw84 & Msm2a4));
	assign Drm2a4 = (Tsm2a4 & Atm2a4);
	assign Atm2a4 = (~(Wsqw84 & Htm2a4));
	assign Tsm2a4 = (~(E6pw84 & Otm2a4));
	assign Pqm2a4 = (Vtm2a4 & Cum2a4);
	assign Cum2a4 = (Jum2a4 & Qum2a4);
	assign Qum2a4 = (~(Ofsw84 & Xum2a4));
	assign Jum2a4 = (~(G2uw84 & Evm2a4));
	assign Vtm2a4 = (Lvm2a4 & Svm2a4);
	assign Svm2a4 = (~(Qbxw84 & Zvm2a4));
	assign Lvm2a4 = (~(Yovw84 & Gwm2a4));
	assign Uim2a4 = (Nwm2a4 | Ltrx84);
	assign Ltrx84 = (!Fizx84);
	assign HWDATA[30] = (~(Uwm2a4 & Bxm2a4));
	assign Bxm2a4 = (Nim2a4 | X41y84);
	assign Uwm2a4 = (Ixm2a4 & Pxm2a4);
	assign Pxm2a4 = (~(N8b2a4 & Dwdx84));
	assign Dwdx84 = (~(Wxm2a4 & Dym2a4));
	assign Dym2a4 = (Kym2a4 & Rym2a4);
	assign Rym2a4 = (Yym2a4 & Fzm2a4);
	assign Fzm2a4 = (Mzm2a4 & Tzm2a4);
	assign Tzm2a4 = (~(Wygw84 & Mlm2a4));
	assign Mzm2a4 = (A0n2a4 & H0n2a4);
	assign H0n2a4 = (~(Ouyw84 & Hmm2a4));
	assign A0n2a4 = (~(Qd0x84 & Omm2a4));
	assign Yym2a4 = (O0n2a4 & V0n2a4);
	assign V0n2a4 = (~(Cgaw84 & Jnm2a4));
	assign O0n2a4 = (~(Oliw84 & Qnm2a4));
	assign Kym2a4 = (C1n2a4 & J1n2a4);
	assign J1n2a4 = (Q1n2a4 & X1n2a4);
	assign X1n2a4 = (~(U2cw84 & Zom2a4));
	assign Q1n2a4 = (~(Mpdw84 & Gpm2a4));
	assign C1n2a4 = (E2n2a4 & L2n2a4);
	assign L2n2a4 = (~(G8kw84 & Bqm2a4));
	assign E2n2a4 = (~(Ecfw84 & Iqm2a4));
	assign Wxm2a4 = (S2n2a4 & Z2n2a4);
	assign Z2n2a4 = (G3n2a4 & N3n2a4);
	assign N3n2a4 = (U3n2a4 & B4n2a4);
	assign B4n2a4 = (~(Yulw84 & Fsm2a4));
	assign U3n2a4 = (~(Qhnw84 & Msm2a4));
	assign G3n2a4 = (I4n2a4 & P4n2a4);
	assign P4n2a4 = (~(Arqw84 & Htm2a4));
	assign I4n2a4 = (~(I4pw84 & Otm2a4));
	assign S2n2a4 = (W4n2a4 & D5n2a4);
	assign D5n2a4 = (K5n2a4 & R5n2a4);
	assign R5n2a4 = (~(Sdsw84 & Xum2a4));
	assign K5n2a4 = (~(K0uw84 & Evm2a4));
	assign W4n2a4 = (Y5n2a4 & F6n2a4);
	assign F6n2a4 = (~(U9xw84 & Zvm2a4));
	assign Y5n2a4 = (~(Cnvw84 & Gwm2a4));
	assign Ixm2a4 = (Nwm2a4 | Akrx84);
	assign HWDATA[2] = (~(Ralx84 | Zhpx84));
	assign HWDATA[29] = (~(M6n2a4 & T6n2a4));
	assign T6n2a4 = (Nim2a4 | Vw0y84);
	assign M6n2a4 = (A7n2a4 & H7n2a4);
	assign H7n2a4 = (~(N8b2a4 & Vitx84));
	assign Vitx84 = (~(O7n2a4 & V7n2a4));
	assign V7n2a4 = (C8n2a4 & J8n2a4);
	assign J8n2a4 = (Q8n2a4 & X8n2a4);
	assign X8n2a4 = (E9n2a4 & L9n2a4);
	assign L9n2a4 = (~(Axgw84 & Mlm2a4));
	assign E9n2a4 = (S9n2a4 & Z9n2a4);
	assign Z9n2a4 = (~(Ssyw84 & Hmm2a4));
	assign S9n2a4 = (~(Ub0x84 & Omm2a4));
	assign Q8n2a4 = (Gan2a4 & Nan2a4);
	assign Nan2a4 = (~(Geaw84 & Jnm2a4));
	assign Gan2a4 = (~(Sjiw84 & Qnm2a4));
	assign C8n2a4 = (Uan2a4 & Bbn2a4);
	assign Bbn2a4 = (Ibn2a4 & Pbn2a4);
	assign Pbn2a4 = (~(Y0cw84 & Zom2a4));
	assign Ibn2a4 = (~(Qndw84 & Gpm2a4));
	assign Uan2a4 = (Wbn2a4 & Dcn2a4);
	assign Dcn2a4 = (~(K6kw84 & Bqm2a4));
	assign Wbn2a4 = (~(Iafw84 & Iqm2a4));
	assign O7n2a4 = (Kcn2a4 & Rcn2a4);
	assign Rcn2a4 = (Ycn2a4 & Fdn2a4);
	assign Fdn2a4 = (Mdn2a4 & Tdn2a4);
	assign Tdn2a4 = (~(Ctlw84 & Fsm2a4));
	assign Mdn2a4 = (~(Ufnw84 & Msm2a4));
	assign Ycn2a4 = (Aen2a4 & Hen2a4);
	assign Hen2a4 = (~(Epqw84 & Htm2a4));
	assign Aen2a4 = (~(M2pw84 & Otm2a4));
	assign Kcn2a4 = (Oen2a4 & Ven2a4);
	assign Ven2a4 = (Cfn2a4 & Jfn2a4);
	assign Jfn2a4 = (~(Wbsw84 & Xum2a4));
	assign Cfn2a4 = (~(Oytw84 & Evm2a4));
	assign Oen2a4 = (Qfn2a4 & Xfn2a4);
	assign Xfn2a4 = (~(Y7xw84 & Zvm2a4));
	assign Qfn2a4 = (~(Glvw84 & Gwm2a4));
	assign A7n2a4 = (Nwm2a4 | Lfrx84);
	assign HWDATA[28] = (~(Egn2a4 & Lgn2a4));
	assign Lgn2a4 = (Nim2a4 | W71y84);
	assign Egn2a4 = (Sgn2a4 & Zgn2a4);
	assign Zgn2a4 = (~(N8b2a4 & W8tx84));
	assign W8tx84 = (~(Ghn2a4 & Nhn2a4));
	assign Nhn2a4 = (Uhn2a4 & Bin2a4);
	assign Bin2a4 = (Iin2a4 & Pin2a4);
	assign Pin2a4 = (Win2a4 & Djn2a4);
	assign Djn2a4 = (~(Evgw84 & Mlm2a4));
	assign Win2a4 = (Kjn2a4 & Rjn2a4);
	assign Rjn2a4 = (~(Wqyw84 & Hmm2a4));
	assign Kjn2a4 = (~(Y90x84 & Omm2a4));
	assign Iin2a4 = (Yjn2a4 & Fkn2a4);
	assign Fkn2a4 = (~(Kcaw84 & Jnm2a4));
	assign Yjn2a4 = (~(Whiw84 & Qnm2a4));
	assign Uhn2a4 = (Mkn2a4 & Tkn2a4);
	assign Tkn2a4 = (Aln2a4 & Hln2a4);
	assign Hln2a4 = (~(Czbw84 & Zom2a4));
	assign Aln2a4 = (~(Uldw84 & Gpm2a4));
	assign Mkn2a4 = (Oln2a4 & Vln2a4);
	assign Vln2a4 = (~(O4kw84 & Bqm2a4));
	assign Oln2a4 = (~(M8fw84 & Iqm2a4));
	assign Ghn2a4 = (Cmn2a4 & Jmn2a4);
	assign Jmn2a4 = (Qmn2a4 & Xmn2a4);
	assign Xmn2a4 = (Enn2a4 & Lnn2a4);
	assign Lnn2a4 = (~(Grlw84 & Fsm2a4));
	assign Enn2a4 = (~(Ydnw84 & Msm2a4));
	assign Qmn2a4 = (Snn2a4 & Znn2a4);
	assign Znn2a4 = (~(Inqw84 & Htm2a4));
	assign Snn2a4 = (~(Q0pw84 & Otm2a4));
	assign Cmn2a4 = (Gon2a4 & Non2a4);
	assign Non2a4 = (Uon2a4 & Bpn2a4);
	assign Bpn2a4 = (~(Aasw84 & Xum2a4));
	assign Uon2a4 = (~(Swtw84 & Evm2a4));
	assign Gon2a4 = (Ipn2a4 & Ppn2a4);
	assign Ppn2a4 = (~(C6xw84 & Zvm2a4));
	assign Ipn2a4 = (~(Kjvw84 & Gwm2a4));
	assign Sgn2a4 = (Nwm2a4 | B01y84);
	assign HWDATA[27] = (~(Wpn2a4 & Dqn2a4));
	assign Dqn2a4 = (Nim2a4 | Tlpx84);
	assign Wpn2a4 = (Kqn2a4 & Rqn2a4);
	assign Rqn2a4 = (Yqn2a4 | E6tx84);
	assign E6tx84 = (Frn2a4 & Mrn2a4);
	assign Mrn2a4 = (Trn2a4 & Asn2a4);
	assign Asn2a4 = (Hsn2a4 & Osn2a4);
	assign Osn2a4 = (Vsn2a4 & Ctn2a4);
	assign Ctn2a4 = (~(Itgw84 & Mlm2a4));
	assign Vsn2a4 = (Jtn2a4 & Qtn2a4);
	assign Qtn2a4 = (~(Apyw84 & Hmm2a4));
	assign Jtn2a4 = (~(C80x84 & Omm2a4));
	assign Hsn2a4 = (Xtn2a4 & Eun2a4);
	assign Eun2a4 = (~(Oaaw84 & Jnm2a4));
	assign Xtn2a4 = (~(Agiw84 & Qnm2a4));
	assign Trn2a4 = (Lun2a4 & Sun2a4);
	assign Sun2a4 = (Zun2a4 & Gvn2a4);
	assign Gvn2a4 = (~(Gxbw84 & Zom2a4));
	assign Zun2a4 = (~(Yjdw84 & Gpm2a4));
	assign Lun2a4 = (Nvn2a4 & Uvn2a4);
	assign Uvn2a4 = (~(S2kw84 & Bqm2a4));
	assign Nvn2a4 = (~(Q6fw84 & Iqm2a4));
	assign Frn2a4 = (Bwn2a4 & Iwn2a4);
	assign Iwn2a4 = (Pwn2a4 & Wwn2a4);
	assign Wwn2a4 = (Dxn2a4 & Kxn2a4);
	assign Kxn2a4 = (~(Kplw84 & Fsm2a4));
	assign Dxn2a4 = (~(Ccnw84 & Msm2a4));
	assign Pwn2a4 = (Rxn2a4 & Yxn2a4);
	assign Yxn2a4 = (~(Mlqw84 & Htm2a4));
	assign Rxn2a4 = (~(Uyow84 & Otm2a4));
	assign Bwn2a4 = (Fyn2a4 & Myn2a4);
	assign Myn2a4 = (Tyn2a4 & Azn2a4);
	assign Azn2a4 = (~(E8sw84 & Xum2a4));
	assign Tyn2a4 = (~(Wutw84 & Evm2a4));
	assign Fyn2a4 = (Hzn2a4 & Ozn2a4);
	assign Ozn2a4 = (~(G4xw84 & Zvm2a4));
	assign Hzn2a4 = (~(Ohvw84 & Gwm2a4));
	assign Kqn2a4 = (Nwm2a4 | H6rx84);
	assign H6rx84 = (!Cdzx84);
	assign HWDATA[26] = (~(Vzn2a4 & C0o2a4));
	assign C0o2a4 = (Nim2a4 | Zhpx84);
	assign Vzn2a4 = (J0o2a4 & Q0o2a4);
	assign Q0o2a4 = (Yqn2a4 | Vxsx84);
	assign Vxsx84 = (!Vczx84);
	assign Vczx84 = (~(X0o2a4 & E1o2a4));
	assign E1o2a4 = (L1o2a4 & S1o2a4);
	assign S1o2a4 = (Z1o2a4 & G2o2a4);
	assign G2o2a4 = (N2o2a4 & U2o2a4);
	assign U2o2a4 = (~(Mrgw84 & Mlm2a4));
	assign N2o2a4 = (B3o2a4 & I3o2a4);
	assign I3o2a4 = (~(Enyw84 & Hmm2a4));
	assign B3o2a4 = (~(G60x84 & Omm2a4));
	assign Z1o2a4 = (P3o2a4 & W3o2a4);
	assign W3o2a4 = (~(S8aw84 & Jnm2a4));
	assign P3o2a4 = (~(Eeiw84 & Qnm2a4));
	assign L1o2a4 = (D4o2a4 & K4o2a4);
	assign K4o2a4 = (R4o2a4 & Y4o2a4);
	assign Y4o2a4 = (~(Kvbw84 & Zom2a4));
	assign R4o2a4 = (~(Cidw84 & Gpm2a4));
	assign D4o2a4 = (F5o2a4 & M5o2a4);
	assign M5o2a4 = (~(W0kw84 & Bqm2a4));
	assign F5o2a4 = (~(U4fw84 & Iqm2a4));
	assign X0o2a4 = (T5o2a4 & A6o2a4);
	assign A6o2a4 = (H6o2a4 & O6o2a4);
	assign O6o2a4 = (V6o2a4 & C7o2a4);
	assign C7o2a4 = (~(Onlw84 & Fsm2a4));
	assign V6o2a4 = (~(Ganw84 & Msm2a4));
	assign H6o2a4 = (J7o2a4 & Q7o2a4);
	assign Q7o2a4 = (~(Qjqw84 & Htm2a4));
	assign J7o2a4 = (~(Ywow84 & Otm2a4));
	assign T5o2a4 = (X7o2a4 & E8o2a4);
	assign E8o2a4 = (L8o2a4 & S8o2a4);
	assign S8o2a4 = (~(I6sw84 & Xum2a4));
	assign L8o2a4 = (~(Attw84 & Evm2a4));
	assign X7o2a4 = (Z8o2a4 & G9o2a4);
	assign G9o2a4 = (~(K2xw84 & Zvm2a4));
	assign Z8o2a4 = (~(Sfvw84 & Gwm2a4));
	assign J0o2a4 = (Nwm2a4 | Yxqx84);
	assign Yxqx84 = (!Sezx84);
	assign HWDATA[25] = (~(N9o2a4 & U9o2a4));
	assign U9o2a4 = (Nim2a4 | Sd0y84);
	assign N9o2a4 = (Bao2a4 & Iao2a4);
	assign Iao2a4 = (Yqn2a4 | Lssx84);
	assign Lssx84 = (!Oczx84);
	assign Oczx84 = (~(Pao2a4 & Wao2a4));
	assign Wao2a4 = (Dbo2a4 & Kbo2a4);
	assign Kbo2a4 = (Rbo2a4 & Ybo2a4);
	assign Ybo2a4 = (Fco2a4 & Mco2a4);
	assign Mco2a4 = (~(Qpgw84 & Mlm2a4));
	assign Fco2a4 = (Tco2a4 & Ado2a4);
	assign Ado2a4 = (~(Ilyw84 & Hmm2a4));
	assign Tco2a4 = (~(K40x84 & Omm2a4));
	assign Rbo2a4 = (Hdo2a4 & Odo2a4);
	assign Odo2a4 = (~(W6aw84 & Jnm2a4));
	assign Hdo2a4 = (~(Iciw84 & Qnm2a4));
	assign Dbo2a4 = (Vdo2a4 & Ceo2a4);
	assign Ceo2a4 = (Jeo2a4 & Qeo2a4);
	assign Qeo2a4 = (~(Otbw84 & Zom2a4));
	assign Jeo2a4 = (~(Ggdw84 & Gpm2a4));
	assign Vdo2a4 = (Xeo2a4 & Efo2a4);
	assign Efo2a4 = (~(Azjw84 & Bqm2a4));
	assign Xeo2a4 = (~(Y2fw84 & Iqm2a4));
	assign Pao2a4 = (Lfo2a4 & Sfo2a4);
	assign Sfo2a4 = (Zfo2a4 & Ggo2a4);
	assign Ggo2a4 = (Ngo2a4 & Ugo2a4);
	assign Ugo2a4 = (~(Sllw84 & Fsm2a4));
	assign Ngo2a4 = (~(K8nw84 & Msm2a4));
	assign Zfo2a4 = (Bho2a4 & Iho2a4);
	assign Iho2a4 = (~(Uhqw84 & Htm2a4));
	assign Bho2a4 = (~(Cvow84 & Otm2a4));
	assign Lfo2a4 = (Pho2a4 & Who2a4);
	assign Who2a4 = (Dio2a4 & Kio2a4);
	assign Kio2a4 = (~(M4sw84 & Xum2a4));
	assign Dio2a4 = (~(Ertw84 & Evm2a4));
	assign Pho2a4 = (Rio2a4 & Yio2a4);
	assign Yio2a4 = (~(O0xw84 & Zvm2a4));
	assign Rio2a4 = (~(Wdvw84 & Gwm2a4));
	assign Bao2a4 = (Nwm2a4 | Cb1y84);
	assign Cb1y84 = (Fjo2a4 & Mjo2a4);
	assign Mjo2a4 = (Tjo2a4 & Ako2a4);
	assign Ako2a4 = (Hko2a4 & Oko2a4);
	assign Oko2a4 = (Vko2a4 & Clo2a4);
	assign Clo2a4 = (~(Dwfw84 & Mlm2a4));
	assign Vko2a4 = (Jlo2a4 & Qlo2a4);
	assign Qlo2a4 = (~(Vrxw84 & Hmm2a4));
	assign Jlo2a4 = (~(Xazw84 & Omm2a4));
	assign Hko2a4 = (Xlo2a4 & Emo2a4);
	assign Emo2a4 = (~(Jd9w84 & Jnm2a4));
	assign Xlo2a4 = (~(Vihw84 & Qnm2a4));
	assign Tjo2a4 = (Lmo2a4 & Smo2a4);
	assign Smo2a4 = (Zmo2a4 & Gno2a4);
	assign Gno2a4 = (~(B0bw84 & Zom2a4));
	assign Zmo2a4 = (~(Tmcw84 & Gpm2a4));
	assign Lmo2a4 = (Nno2a4 & Uno2a4);
	assign Uno2a4 = (~(N5jw84 & Bqm2a4));
	assign Nno2a4 = (~(L9ew84 & Iqm2a4));
	assign Fjo2a4 = (Boo2a4 & Ioo2a4);
	assign Ioo2a4 = (Poo2a4 & Woo2a4);
	assign Woo2a4 = (Dpo2a4 & Kpo2a4);
	assign Kpo2a4 = (~(Fskw84 & Fsm2a4));
	assign Dpo2a4 = (~(Xemw84 & Msm2a4));
	assign Poo2a4 = (Rpo2a4 & Ypo2a4);
	assign Ypo2a4 = (~(Hopw84 & Htm2a4));
	assign Rpo2a4 = (~(P1ow84 & Otm2a4));
	assign Boo2a4 = (Fqo2a4 & Mqo2a4);
	assign Mqo2a4 = (Tqo2a4 & Aro2a4);
	assign Aro2a4 = (~(Zarw84 & Xum2a4));
	assign Tqo2a4 = (~(Rxsw84 & Evm2a4));
	assign Fqo2a4 = (Hro2a4 & Oro2a4);
	assign Oro2a4 = (~(B7ww84 & Zvm2a4));
	assign Hro2a4 = (~(Jkuw84 & Gwm2a4));
	assign HWDATA[24] = (~(Vro2a4 & Cso2a4));
	assign Cso2a4 = (Nim2a4 | Yn0y84);
	assign Vro2a4 = (Jso2a4 & Qso2a4);
	assign Qso2a4 = (Nwm2a4 | M21y84);
	assign M21y84 = (Xso2a4 & Eto2a4);
	assign Eto2a4 = (Lto2a4 & Sto2a4);
	assign Sto2a4 = (Zto2a4 & Guo2a4);
	assign Guo2a4 = (Nuo2a4 & Uuo2a4);
	assign Uuo2a4 = (~(Iufw84 & Mlm2a4));
	assign Nuo2a4 = (Bvo2a4 & Ivo2a4);
	assign Ivo2a4 = (~(Aqxw84 & Hmm2a4));
	assign Bvo2a4 = (~(C9zw84 & Omm2a4));
	assign Zto2a4 = (Pvo2a4 & Wvo2a4);
	assign Wvo2a4 = (~(Ob9w84 & Jnm2a4));
	assign Pvo2a4 = (~(Ahhw84 & Qnm2a4));
	assign Lto2a4 = (Dwo2a4 & Kwo2a4);
	assign Kwo2a4 = (Rwo2a4 & Ywo2a4);
	assign Ywo2a4 = (~(Gyaw84 & Zom2a4));
	assign Rwo2a4 = (~(Ykcw84 & Gpm2a4));
	assign Dwo2a4 = (Fxo2a4 & Mxo2a4);
	assign Mxo2a4 = (~(S3jw84 & Bqm2a4));
	assign Fxo2a4 = (~(Q7ew84 & Iqm2a4));
	assign Xso2a4 = (Txo2a4 & Ayo2a4);
	assign Ayo2a4 = (Hyo2a4 & Oyo2a4);
	assign Oyo2a4 = (Vyo2a4 & Czo2a4);
	assign Czo2a4 = (~(Kqkw84 & Fsm2a4));
	assign Vyo2a4 = (~(Cdmw84 & Msm2a4));
	assign Hyo2a4 = (Jzo2a4 & Qzo2a4);
	assign Qzo2a4 = (~(Mmpw84 & Htm2a4));
	assign Jzo2a4 = (~(Uznw84 & Otm2a4));
	assign Txo2a4 = (Xzo2a4 & E0p2a4);
	assign E0p2a4 = (L0p2a4 & S0p2a4);
	assign S0p2a4 = (~(E9rw84 & Xum2a4));
	assign L0p2a4 = (~(Wvsw84 & Evm2a4));
	assign Xzo2a4 = (Z0p2a4 & G1p2a4);
	assign G1p2a4 = (~(G5ww84 & Zvm2a4));
	assign Z0p2a4 = (~(Oiuw84 & Gwm2a4));
	assign Nwm2a4 = (N1p2a4 | Ralx84);
	assign Jso2a4 = (Yqn2a4 | Yf1y84);
	assign Yf1y84 = (U1p2a4 & B2p2a4);
	assign B2p2a4 = (I2p2a4 & P2p2a4);
	assign P2p2a4 = (W2p2a4 & D3p2a4);
	assign D3p2a4 = (K3p2a4 & R3p2a4);
	assign R3p2a4 = (~(Ungw84 & Mlm2a4));
	assign K3p2a4 = (Y3p2a4 & F4p2a4);
	assign F4p2a4 = (~(Mjyw84 & Hmm2a4));
	assign Y3p2a4 = (~(O20x84 & Omm2a4));
	assign W2p2a4 = (M4p2a4 & T4p2a4);
	assign T4p2a4 = (~(A5aw84 & Jnm2a4));
	assign M4p2a4 = (~(Maiw84 & Qnm2a4));
	assign I2p2a4 = (A5p2a4 & H5p2a4);
	assign H5p2a4 = (O5p2a4 & V5p2a4);
	assign V5p2a4 = (~(Srbw84 & Zom2a4));
	assign O5p2a4 = (~(Kedw84 & Gpm2a4));
	assign A5p2a4 = (C6p2a4 & J6p2a4);
	assign J6p2a4 = (~(Exjw84 & Bqm2a4));
	assign C6p2a4 = (~(C1fw84 & Iqm2a4));
	assign U1p2a4 = (Q6p2a4 & X6p2a4);
	assign X6p2a4 = (E7p2a4 & L7p2a4);
	assign L7p2a4 = (S7p2a4 & Z7p2a4);
	assign Z7p2a4 = (~(Wjlw84 & Fsm2a4));
	assign S7p2a4 = (~(O6nw84 & Msm2a4));
	assign E7p2a4 = (G8p2a4 & N8p2a4);
	assign N8p2a4 = (~(Yfqw84 & Htm2a4));
	assign G8p2a4 = (~(Gtow84 & Otm2a4));
	assign Q6p2a4 = (U8p2a4 & B9p2a4);
	assign B9p2a4 = (I9p2a4 & P9p2a4);
	assign P9p2a4 = (~(Q2sw84 & Xum2a4));
	assign I9p2a4 = (~(Iptw84 & Evm2a4));
	assign U8p2a4 = (W9p2a4 & Dap2a4);
	assign Dap2a4 = (~(Syww84 & Zvm2a4));
	assign W9p2a4 = (~(Acvw84 & Gwm2a4));
	assign HWDATA[23] = (!Ezex84);
	assign Ezex84 = (N8b2a4 ? Xksx84 : Piqx84);
	assign Xksx84 = (!Lezx84);
	assign Lezx84 = (~(Kap2a4 & Rap2a4));
	assign Rap2a4 = (Yap2a4 & Fbp2a4);
	assign Fbp2a4 = (Mbp2a4 & Tbp2a4);
	assign Tbp2a4 = (Acp2a4 & Hcp2a4);
	assign Hcp2a4 = (~(Ylgw84 & Mlm2a4));
	assign Acp2a4 = (Ocp2a4 & Vcp2a4);
	assign Vcp2a4 = (~(Qhyw84 & Hmm2a4));
	assign Ocp2a4 = (~(S00x84 & Omm2a4));
	assign Mbp2a4 = (Cdp2a4 & Jdp2a4);
	assign Jdp2a4 = (~(E3aw84 & Jnm2a4));
	assign Cdp2a4 = (~(Q8iw84 & Qnm2a4));
	assign Yap2a4 = (Qdp2a4 & Xdp2a4);
	assign Xdp2a4 = (Eep2a4 & Lep2a4);
	assign Lep2a4 = (~(Wpbw84 & Zom2a4));
	assign Eep2a4 = (~(Ocdw84 & Gpm2a4));
	assign Qdp2a4 = (Sep2a4 & Zep2a4);
	assign Zep2a4 = (~(Ivjw84 & Bqm2a4));
	assign Sep2a4 = (~(Gzew84 & Iqm2a4));
	assign Kap2a4 = (Gfp2a4 & Nfp2a4);
	assign Nfp2a4 = (Ufp2a4 & Bgp2a4);
	assign Bgp2a4 = (Igp2a4 & Pgp2a4);
	assign Pgp2a4 = (~(Ailw84 & Fsm2a4));
	assign Igp2a4 = (~(S4nw84 & Msm2a4));
	assign Ufp2a4 = (Wgp2a4 & Dhp2a4);
	assign Dhp2a4 = (~(Ceqw84 & Htm2a4));
	assign Wgp2a4 = (~(Krow84 & Otm2a4));
	assign Gfp2a4 = (Khp2a4 & Rhp2a4);
	assign Rhp2a4 = (Yhp2a4 & Fip2a4);
	assign Fip2a4 = (~(U0sw84 & Xum2a4));
	assign Yhp2a4 = (~(Mntw84 & Evm2a4));
	assign Khp2a4 = (Mip2a4 & Tip2a4);
	assign Tip2a4 = (~(Wwww84 & Zvm2a4));
	assign Mip2a4 = (~(Eavw84 & Gwm2a4));
	assign Piqx84 = (!Mizx84);
	assign HWDATA[22] = (!Ajp2a4);
	assign Ajp2a4 = (N8b2a4 ? Fisx84 : X41y84);
	assign Fisx84 = (!Igzx84);
	assign Igzx84 = (~(Hjp2a4 & Ojp2a4));
	assign Ojp2a4 = (Vjp2a4 & Ckp2a4);
	assign Ckp2a4 = (Jkp2a4 & Qkp2a4);
	assign Qkp2a4 = (Xkp2a4 & Elp2a4);
	assign Elp2a4 = (~(Ckgw84 & Mlm2a4));
	assign Xkp2a4 = (Llp2a4 & Slp2a4);
	assign Slp2a4 = (~(Ufyw84 & Hmm2a4));
	assign Llp2a4 = (~(Wyzw84 & Omm2a4));
	assign Jkp2a4 = (Zlp2a4 & Gmp2a4);
	assign Gmp2a4 = (~(I1aw84 & Jnm2a4));
	assign Zlp2a4 = (~(U6iw84 & Qnm2a4));
	assign Vjp2a4 = (Nmp2a4 & Ump2a4);
	assign Ump2a4 = (Bnp2a4 & Inp2a4);
	assign Inp2a4 = (~(Aobw84 & Zom2a4));
	assign Bnp2a4 = (~(Sadw84 & Gpm2a4));
	assign Nmp2a4 = (Pnp2a4 & Wnp2a4);
	assign Wnp2a4 = (~(Mtjw84 & Bqm2a4));
	assign Pnp2a4 = (~(Kxew84 & Iqm2a4));
	assign Hjp2a4 = (Dop2a4 & Kop2a4);
	assign Kop2a4 = (Rop2a4 & Yop2a4);
	assign Yop2a4 = (Fpp2a4 & Mpp2a4);
	assign Mpp2a4 = (~(Eglw84 & Fsm2a4));
	assign Fpp2a4 = (~(W2nw84 & Msm2a4));
	assign Rop2a4 = (Tpp2a4 & Aqp2a4);
	assign Aqp2a4 = (~(Gcqw84 & Htm2a4));
	assign Tpp2a4 = (~(Opow84 & Otm2a4));
	assign Dop2a4 = (Hqp2a4 & Oqp2a4);
	assign Oqp2a4 = (Vqp2a4 & Crp2a4);
	assign Crp2a4 = (~(Yyrw84 & Xum2a4));
	assign Vqp2a4 = (~(Qltw84 & Evm2a4));
	assign Hqp2a4 = (Jrp2a4 & Qrp2a4);
	assign Qrp2a4 = (~(Avww84 & Zvm2a4));
	assign Jrp2a4 = (~(I8vw84 & Gwm2a4));
	assign HWDATA[21] = (!Z7b2a4);
	assign Z7b2a4 = (N8b2a4 ? Qdsx84 : Vw0y84);
	assign Qdsx84 = (!Wgzx84);
	assign Wgzx84 = (~(Xrp2a4 & Esp2a4));
	assign Esp2a4 = (Lsp2a4 & Ssp2a4);
	assign Ssp2a4 = (Zsp2a4 & Gtp2a4);
	assign Gtp2a4 = (Ntp2a4 & Utp2a4);
	assign Utp2a4 = (~(Gigw84 & Mlm2a4));
	assign Ntp2a4 = (Bup2a4 & Iup2a4);
	assign Iup2a4 = (~(Ydyw84 & Hmm2a4));
	assign Bup2a4 = (~(Axzw84 & Omm2a4));
	assign Zsp2a4 = (Pup2a4 & Wup2a4);
	assign Wup2a4 = (~(Mz9w84 & Jnm2a4));
	assign Pup2a4 = (~(Y4iw84 & Qnm2a4));
	assign Lsp2a4 = (Dvp2a4 & Kvp2a4);
	assign Kvp2a4 = (Rvp2a4 & Yvp2a4);
	assign Yvp2a4 = (~(Embw84 & Zom2a4));
	assign Rvp2a4 = (~(W8dw84 & Gpm2a4));
	assign Dvp2a4 = (Fwp2a4 & Mwp2a4);
	assign Mwp2a4 = (~(Qrjw84 & Bqm2a4));
	assign Fwp2a4 = (~(Ovew84 & Iqm2a4));
	assign Xrp2a4 = (Twp2a4 & Axp2a4);
	assign Axp2a4 = (Hxp2a4 & Oxp2a4);
	assign Oxp2a4 = (Vxp2a4 & Cyp2a4);
	assign Cyp2a4 = (~(Ielw84 & Fsm2a4));
	assign Vxp2a4 = (~(A1nw84 & Msm2a4));
	assign Hxp2a4 = (Jyp2a4 & Qyp2a4);
	assign Qyp2a4 = (~(Kaqw84 & Htm2a4));
	assign Jyp2a4 = (~(Snow84 & Otm2a4));
	assign Twp2a4 = (Xyp2a4 & Ezp2a4);
	assign Ezp2a4 = (Lzp2a4 & Szp2a4);
	assign Szp2a4 = (~(Cxrw84 & Xum2a4));
	assign Lzp2a4 = (~(Ujtw84 & Evm2a4));
	assign Xyp2a4 = (Zzp2a4 & G0q2a4);
	assign G0q2a4 = (~(Etww84 & Zvm2a4));
	assign Zzp2a4 = (~(M6vw84 & Gwm2a4));
	assign HWDATA[20] = (Yqn2a4 ? Shm2a4 : Pgzx84);
	assign Yqn2a4 = (!N8b2a4);
	assign Pgzx84 = (~(N0q2a4 & U0q2a4));
	assign U0q2a4 = (B1q2a4 & I1q2a4);
	assign I1q2a4 = (P1q2a4 & W1q2a4);
	assign W1q2a4 = (D2q2a4 & K2q2a4);
	assign K2q2a4 = (~(Kggw84 & Mlm2a4));
	assign D2q2a4 = (R2q2a4 & Y2q2a4);
	assign Y2q2a4 = (~(Ccyw84 & Hmm2a4));
	assign R2q2a4 = (~(Evzw84 & Omm2a4));
	assign P1q2a4 = (F3q2a4 & M3q2a4);
	assign M3q2a4 = (~(Qx9w84 & Jnm2a4));
	assign F3q2a4 = (~(C3iw84 & Qnm2a4));
	assign B1q2a4 = (T3q2a4 & A4q2a4);
	assign A4q2a4 = (H4q2a4 & O4q2a4);
	assign O4q2a4 = (~(Ikbw84 & Zom2a4));
	assign H4q2a4 = (~(A7dw84 & Gpm2a4));
	assign T3q2a4 = (V4q2a4 & C5q2a4);
	assign C5q2a4 = (~(Upjw84 & Bqm2a4));
	assign V4q2a4 = (~(Stew84 & Iqm2a4));
	assign N0q2a4 = (J5q2a4 & Q5q2a4);
	assign Q5q2a4 = (X5q2a4 & E6q2a4);
	assign E6q2a4 = (L6q2a4 & S6q2a4);
	assign S6q2a4 = (~(Mclw84 & Fsm2a4));
	assign L6q2a4 = (~(Ezmw84 & Msm2a4));
	assign X5q2a4 = (Z6q2a4 & G7q2a4);
	assign G7q2a4 = (~(O8qw84 & Htm2a4));
	assign Z6q2a4 = (~(Wlow84 & Otm2a4));
	assign J5q2a4 = (N7q2a4 & U7q2a4);
	assign U7q2a4 = (B8q2a4 & I8q2a4);
	assign I8q2a4 = (~(Gvrw84 & Xum2a4));
	assign B8q2a4 = (~(Yhtw84 & Evm2a4));
	assign N7q2a4 = (P8q2a4 & W8q2a4);
	assign W8q2a4 = (~(Irww84 & Zvm2a4));
	assign P8q2a4 = (~(Q4vw84 & Gwm2a4));
	assign HWDATA[1] = (~(Ralx84 | Sd0y84));
	assign HWDATA[19] = (!S7b2a4);
	assign S7b2a4 = (N8b2a4 ? Du0y84 : Tlpx84);
	assign Du0y84 = (D9q2a4 & K9q2a4);
	assign K9q2a4 = (R9q2a4 & Y9q2a4);
	assign Y9q2a4 = (Faq2a4 & Maq2a4);
	assign Maq2a4 = (Taq2a4 & Abq2a4);
	assign Abq2a4 = (~(Oegw84 & Mlm2a4));
	assign Taq2a4 = (Hbq2a4 & Obq2a4);
	assign Obq2a4 = (~(Gayw84 & Hmm2a4));
	assign Hbq2a4 = (~(Itzw84 & Omm2a4));
	assign Faq2a4 = (Vbq2a4 & Ccq2a4);
	assign Ccq2a4 = (~(Uv9w84 & Jnm2a4));
	assign Vbq2a4 = (~(G1iw84 & Qnm2a4));
	assign R9q2a4 = (Jcq2a4 & Qcq2a4);
	assign Qcq2a4 = (Xcq2a4 & Edq2a4);
	assign Edq2a4 = (~(Mibw84 & Zom2a4));
	assign Xcq2a4 = (~(E5dw84 & Gpm2a4));
	assign Jcq2a4 = (Ldq2a4 & Sdq2a4);
	assign Sdq2a4 = (~(Ynjw84 & Bqm2a4));
	assign Ldq2a4 = (~(Wrew84 & Iqm2a4));
	assign D9q2a4 = (Zdq2a4 & Geq2a4);
	assign Geq2a4 = (Neq2a4 & Ueq2a4);
	assign Ueq2a4 = (Bfq2a4 & Ifq2a4);
	assign Ifq2a4 = (~(Qalw84 & Fsm2a4));
	assign Bfq2a4 = (~(Ixmw84 & Msm2a4));
	assign Neq2a4 = (Pfq2a4 & Wfq2a4);
	assign Wfq2a4 = (~(S6qw84 & Htm2a4));
	assign Pfq2a4 = (~(Akow84 & Otm2a4));
	assign Zdq2a4 = (Dgq2a4 & Kgq2a4);
	assign Kgq2a4 = (Rgq2a4 & Ygq2a4);
	assign Ygq2a4 = (~(Ktrw84 & Xum2a4));
	assign Rgq2a4 = (~(Cgtw84 & Evm2a4));
	assign Dgq2a4 = (Fhq2a4 & Mhq2a4);
	assign Mhq2a4 = (~(Mpww84 & Zvm2a4));
	assign Fhq2a4 = (~(U2vw84 & Gwm2a4));
	assign Tlpx84 = (!Yhzx84);
	assign HWDATA[18] = (!Thq2a4);
	assign Thq2a4 = (N8b2a4 ? Sr0y84 : Zhpx84);
	assign Sr0y84 = (Aiq2a4 & Hiq2a4);
	assign Hiq2a4 = (Oiq2a4 & Viq2a4);
	assign Viq2a4 = (Cjq2a4 & Jjq2a4);
	assign Jjq2a4 = (Qjq2a4 & Xjq2a4);
	assign Xjq2a4 = (~(Scgw84 & Mlm2a4));
	assign Qjq2a4 = (Ekq2a4 & Lkq2a4);
	assign Lkq2a4 = (~(K8yw84 & Hmm2a4));
	assign Ekq2a4 = (~(Mrzw84 & Omm2a4));
	assign Cjq2a4 = (Skq2a4 & Zkq2a4);
	assign Zkq2a4 = (~(Yt9w84 & Jnm2a4));
	assign Skq2a4 = (~(Kzhw84 & Qnm2a4));
	assign Oiq2a4 = (Glq2a4 & Nlq2a4);
	assign Nlq2a4 = (Ulq2a4 & Bmq2a4);
	assign Bmq2a4 = (~(Qgbw84 & Zom2a4));
	assign Ulq2a4 = (~(I3dw84 & Gpm2a4));
	assign Glq2a4 = (Imq2a4 & Pmq2a4);
	assign Pmq2a4 = (~(Cmjw84 & Bqm2a4));
	assign Imq2a4 = (~(Aqew84 & Iqm2a4));
	assign Aiq2a4 = (Wmq2a4 & Dnq2a4);
	assign Dnq2a4 = (Knq2a4 & Rnq2a4);
	assign Rnq2a4 = (Ynq2a4 & Foq2a4);
	assign Foq2a4 = (~(U8lw84 & Fsm2a4));
	assign Ynq2a4 = (~(Mvmw84 & Msm2a4));
	assign Knq2a4 = (Moq2a4 & Toq2a4);
	assign Toq2a4 = (~(W4qw84 & Htm2a4));
	assign Moq2a4 = (~(Eiow84 & Otm2a4));
	assign Wmq2a4 = (Apq2a4 & Hpq2a4);
	assign Hpq2a4 = (Opq2a4 & Vpq2a4);
	assign Vpq2a4 = (~(Orrw84 & Xum2a4));
	assign Opq2a4 = (~(Getw84 & Evm2a4));
	assign Apq2a4 = (Cqq2a4 & Jqq2a4);
	assign Jqq2a4 = (~(Qnww84 & Zvm2a4));
	assign Cqq2a4 = (~(Y0vw84 & Gwm2a4));
	assign Zhpx84 = (!Rhzx84);
	assign HWDATA[17] = (!C6b2a4);
	assign C6b2a4 = (N8b2a4 ? Nd1y84 : Sd0y84);
	assign Nd1y84 = (Qqq2a4 & Xqq2a4);
	assign Xqq2a4 = (Erq2a4 & Lrq2a4);
	assign Lrq2a4 = (Srq2a4 & Zrq2a4);
	assign Zrq2a4 = (Gsq2a4 & Nsq2a4);
	assign Nsq2a4 = (~(Wagw84 & Mlm2a4));
	assign Gsq2a4 = (Usq2a4 & Btq2a4);
	assign Btq2a4 = (~(O6yw84 & Hmm2a4));
	assign Usq2a4 = (~(Qpzw84 & Omm2a4));
	assign Srq2a4 = (Itq2a4 & Ptq2a4);
	assign Ptq2a4 = (~(Cs9w84 & Jnm2a4));
	assign Itq2a4 = (~(Oxhw84 & Qnm2a4));
	assign Erq2a4 = (Wtq2a4 & Duq2a4);
	assign Duq2a4 = (Kuq2a4 & Ruq2a4);
	assign Ruq2a4 = (~(Uebw84 & Zom2a4));
	assign Kuq2a4 = (~(M1dw84 & Gpm2a4));
	assign Wtq2a4 = (Yuq2a4 & Fvq2a4);
	assign Fvq2a4 = (~(Gkjw84 & Bqm2a4));
	assign Yuq2a4 = (~(Eoew84 & Iqm2a4));
	assign Qqq2a4 = (Mvq2a4 & Tvq2a4);
	assign Tvq2a4 = (Awq2a4 & Hwq2a4);
	assign Hwq2a4 = (Owq2a4 & Vwq2a4);
	assign Vwq2a4 = (~(Y6lw84 & Fsm2a4));
	assign Owq2a4 = (~(Qtmw84 & Msm2a4));
	assign Awq2a4 = (Cxq2a4 & Jxq2a4);
	assign Jxq2a4 = (~(A3qw84 & Htm2a4));
	assign Cxq2a4 = (~(Igow84 & Otm2a4));
	assign Mvq2a4 = (Qxq2a4 & Xxq2a4);
	assign Xxq2a4 = (Eyq2a4 & Lyq2a4);
	assign Lyq2a4 = (~(Sprw84 & Xum2a4));
	assign Eyq2a4 = (~(Kctw84 & Evm2a4));
	assign Qxq2a4 = (Syq2a4 & Zyq2a4);
	assign Zyq2a4 = (~(Ulww84 & Zvm2a4));
	assign Syq2a4 = (~(Czuw84 & Gwm2a4));
	assign Sd0y84 = (!Y8gx84);
	assign Y8gx84 = (~(Gzq2a4 & Nzq2a4));
	assign Nzq2a4 = (Uzq2a4 & B0r2a4);
	assign B0r2a4 = (I0r2a4 & P0r2a4);
	assign P0r2a4 = (~(Rhfw84 & Mlm2a4));
	assign I0r2a4 = (~(Xy8w84 & Jnm2a4));
	assign Uzq2a4 = (W0r2a4 & D1r2a4);
	assign D1r2a4 = (~(J4hw84 & Qnm2a4));
	assign W0r2a4 = (~(Plaw84 & Zom2a4));
	assign Gzq2a4 = (K1r2a4 & R1r2a4);
	assign R1r2a4 = (Y1r2a4 & F2r2a4);
	assign F2r2a4 = (~(H8cw84 & Gpm2a4));
	assign Y1r2a4 = (~(Briw84 & Bqm2a4));
	assign K1r2a4 = (Rmk2a4 & M2r2a4);
	assign M2r2a4 = (~(Zudw84 & Iqm2a4));
	assign Rmk2a4 = (T2r2a4 & A3r2a4);
	assign A3r2a4 = (H3r2a4 & O3r2a4);
	assign O3r2a4 = (V3r2a4 & C4r2a4);
	assign C4r2a4 = (~(Fjsw84 & Evm2a4));
	assign V3r2a4 = (~(L0mw84 & Msm2a4));
	assign H3r2a4 = (J4r2a4 & Q4r2a4);
	assign Q4r2a4 = (~(Dnnw84 & Otm2a4));
	assign J4r2a4 = (~(V9pw84 & Htm2a4));
	assign T2r2a4 = (X4r2a4 & E5r2a4);
	assign E5r2a4 = (L5r2a4 & S5r2a4);
	assign S5r2a4 = (~(X5uw84 & Gwm2a4));
	assign L5r2a4 = (~(Psvw84 & Zvm2a4));
	assign X4r2a4 = (Z5r2a4 & G6r2a4);
	assign G6r2a4 = (~(Nwqw84 & Xum2a4));
	assign Z5r2a4 = (~(Tdkw84 & Fsm2a4));
	assign HWDATA[16] = (!W1fx84);
	assign W1fx84 = (N8b2a4 ? Vhux84 : Yn0y84);
	assign N8b2a4 = (~(Ralx84 | N6r2a4));
	assign Vhux84 = (!Bgzx84);
	assign Bgzx84 = (~(U6r2a4 & B7r2a4));
	assign B7r2a4 = (I7r2a4 & P7r2a4);
	assign P7r2a4 = (W7r2a4 & D8r2a4);
	assign D8r2a4 = (K8r2a4 & R8r2a4);
	assign R8r2a4 = (~(A9gw84 & Mlm2a4));
	assign K8r2a4 = (Y8r2a4 & F9r2a4);
	assign F9r2a4 = (~(S4yw84 & Hmm2a4));
	assign Y8r2a4 = (~(Unzw84 & Omm2a4));
	assign W7r2a4 = (M9r2a4 & T9r2a4);
	assign T9r2a4 = (~(Gq9w84 & Jnm2a4));
	assign M9r2a4 = (~(Svhw84 & Qnm2a4));
	assign I7r2a4 = (Aar2a4 & Har2a4);
	assign Har2a4 = (Oar2a4 & Var2a4);
	assign Var2a4 = (~(Ycbw84 & Zom2a4));
	assign Oar2a4 = (~(Qzcw84 & Gpm2a4));
	assign Aar2a4 = (Cbr2a4 & Jbr2a4);
	assign Jbr2a4 = (~(Kijw84 & Bqm2a4));
	assign Cbr2a4 = (~(Imew84 & Iqm2a4));
	assign U6r2a4 = (Qbr2a4 & Xbr2a4);
	assign Xbr2a4 = (Ecr2a4 & Lcr2a4);
	assign Lcr2a4 = (Scr2a4 & Zcr2a4);
	assign Zcr2a4 = (~(C5lw84 & Fsm2a4));
	assign Scr2a4 = (~(Urmw84 & Msm2a4));
	assign Ecr2a4 = (Gdr2a4 & Ndr2a4);
	assign Ndr2a4 = (~(E1qw84 & Htm2a4));
	assign Gdr2a4 = (~(Meow84 & Otm2a4));
	assign Qbr2a4 = (Udr2a4 & Ber2a4);
	assign Ber2a4 = (Ier2a4 & Per2a4);
	assign Per2a4 = (~(Wnrw84 & Xum2a4));
	assign Ier2a4 = (~(Oatw84 & Evm2a4));
	assign Udr2a4 = (Wer2a4 & Dfr2a4);
	assign Dfr2a4 = (~(Yjww84 & Zvm2a4));
	assign Wer2a4 = (~(Gxuw84 & Gwm2a4));
	assign HWDATA[15] = (Nim2a4 ? Fizx84 : Mizx84);
	assign Fizx84 = (~(Kfr2a4 & Rfr2a4));
	assign Rfr2a4 = (Yfr2a4 & Fgr2a4);
	assign Fgr2a4 = (Mgr2a4 & Tgr2a4);
	assign Tgr2a4 = (Ahr2a4 & Hhr2a4);
	assign Hhr2a4 = (~(E7gw84 & Mlm2a4));
	assign Ahr2a4 = (Ohr2a4 & Vhr2a4);
	assign Vhr2a4 = (~(W2yw84 & Hmm2a4));
	assign Ohr2a4 = (~(Ylzw84 & Omm2a4));
	assign Mgr2a4 = (Cir2a4 & Jir2a4);
	assign Jir2a4 = (~(Ko9w84 & Jnm2a4));
	assign Cir2a4 = (~(Wthw84 & Qnm2a4));
	assign Yfr2a4 = (Qir2a4 & Xir2a4);
	assign Xir2a4 = (Ejr2a4 & Ljr2a4);
	assign Ljr2a4 = (~(Cbbw84 & Zom2a4));
	assign Ejr2a4 = (~(Uxcw84 & Gpm2a4));
	assign Qir2a4 = (Sjr2a4 & Zjr2a4);
	assign Zjr2a4 = (~(Ogjw84 & Bqm2a4));
	assign Sjr2a4 = (~(Mkew84 & Iqm2a4));
	assign Kfr2a4 = (Gkr2a4 & Nkr2a4);
	assign Nkr2a4 = (Ukr2a4 & Blr2a4);
	assign Blr2a4 = (Ilr2a4 & Plr2a4);
	assign Plr2a4 = (~(G3lw84 & Fsm2a4));
	assign Ilr2a4 = (~(Ypmw84 & Msm2a4));
	assign Ukr2a4 = (Wlr2a4 & Dmr2a4);
	assign Dmr2a4 = (~(Izpw84 & Htm2a4));
	assign Wlr2a4 = (~(Qcow84 & Otm2a4));
	assign Gkr2a4 = (Kmr2a4 & Rmr2a4);
	assign Rmr2a4 = (Ymr2a4 & Fnr2a4);
	assign Fnr2a4 = (~(Amrw84 & Xum2a4));
	assign Ymr2a4 = (~(S8tw84 & Evm2a4));
	assign Kmr2a4 = (Mnr2a4 & Tnr2a4);
	assign Tnr2a4 = (~(Ciww84 & Zvm2a4));
	assign Mnr2a4 = (~(Kvuw84 & Gwm2a4));
	assign Mizx84 = (~(Aor2a4 & Hor2a4));
	assign Hor2a4 = (Oor2a4 & Vor2a4);
	assign Vor2a4 = (Cpr2a4 & Jpr2a4);
	assign Jpr2a4 = (~(Nsfw84 & Mlm2a4));
	assign Cpr2a4 = (Qpr2a4 & Xpr2a4);
	assign Xpr2a4 = (~(Foxw84 & Hmm2a4));
	assign Qpr2a4 = (~(H7zw84 & Omm2a4));
	assign Oor2a4 = (Eqr2a4 & Lqr2a4);
	assign Lqr2a4 = (~(T99w84 & Jnm2a4));
	assign Eqr2a4 = (~(Ffhw84 & Qnm2a4));
	assign Aor2a4 = (Sqr2a4 & Zqr2a4);
	assign Zqr2a4 = (Grr2a4 & Nrr2a4);
	assign Nrr2a4 = (~(X1jw84 & Bqm2a4));
	assign Grr2a4 = (Urr2a4 & Bsr2a4);
	assign Bsr2a4 = (~(Lwaw84 & Zom2a4));
	assign Urr2a4 = (~(Djcw84 & Gpm2a4));
	assign Sqr2a4 = (Vhk2a4 & Isr2a4);
	assign Isr2a4 = (~(V5ew84 & Iqm2a4));
	assign Vhk2a4 = (Psr2a4 & Wsr2a4);
	assign Wsr2a4 = (Dtr2a4 & Ktr2a4);
	assign Ktr2a4 = (Rtr2a4 & Ytr2a4);
	assign Ytr2a4 = (~(L3ww84 & Zvm2a4));
	assign Rtr2a4 = (~(Busw84 & Evm2a4));
	assign Dtr2a4 = (Fur2a4 & Mur2a4);
	assign Mur2a4 = (~(Zxnw84 & Otm2a4));
	assign Fur2a4 = (~(Rkpw84 & Htm2a4));
	assign Psr2a4 = (Tur2a4 & Avr2a4);
	assign Avr2a4 = (Hvr2a4 & Ovr2a4);
	assign Ovr2a4 = (~(Pokw84 & Fsm2a4));
	assign Hvr2a4 = (~(J7rw84 & Xum2a4));
	assign Tur2a4 = (Vvr2a4 & Cwr2a4);
	assign Cwr2a4 = (~(Tguw84 & Gwm2a4));
	assign Vvr2a4 = (~(Hbmw84 & Msm2a4));
	assign HWDATA[14] = (!Jwr2a4);
	assign Jwr2a4 = (Ehm2a4 ? X41y84 : Akrx84);
	assign X41y84 = (Qwr2a4 & Xwr2a4);
	assign Xwr2a4 = (Exr2a4 & Lxr2a4);
	assign Lxr2a4 = (Sxr2a4 & Zxr2a4);
	assign Zxr2a4 = (~(Sqfw84 & Mlm2a4));
	assign Sxr2a4 = (Gyr2a4 & Nyr2a4);
	assign Nyr2a4 = (~(Kmxw84 & Hmm2a4));
	assign Gyr2a4 = (~(M5zw84 & Omm2a4));
	assign Exr2a4 = (Uyr2a4 & Bzr2a4);
	assign Bzr2a4 = (~(Y79w84 & Jnm2a4));
	assign Uyr2a4 = (~(Kdhw84 & Qnm2a4));
	assign Qwr2a4 = (Izr2a4 & Pzr2a4);
	assign Pzr2a4 = (Wzr2a4 & D0s2a4);
	assign D0s2a4 = (~(C0jw84 & Bqm2a4));
	assign Wzr2a4 = (K0s2a4 & R0s2a4);
	assign R0s2a4 = (~(Quaw84 & Zom2a4));
	assign K0s2a4 = (~(Ihcw84 & Gpm2a4));
	assign Izr2a4 = (Ohk2a4 & Y0s2a4);
	assign Y0s2a4 = (~(A4ew84 & Iqm2a4));
	assign Ohk2a4 = (F1s2a4 & M1s2a4);
	assign M1s2a4 = (T1s2a4 & A2s2a4);
	assign A2s2a4 = (H2s2a4 & O2s2a4);
	assign O2s2a4 = (~(Q1ww84 & Zvm2a4));
	assign H2s2a4 = (~(Gssw84 & Evm2a4));
	assign T1s2a4 = (V2s2a4 & C3s2a4);
	assign C3s2a4 = (~(Ewnw84 & Otm2a4));
	assign V2s2a4 = (~(Wipw84 & Htm2a4));
	assign F1s2a4 = (J3s2a4 & Q3s2a4);
	assign Q3s2a4 = (X3s2a4 & E4s2a4);
	assign E4s2a4 = (~(Umkw84 & Fsm2a4));
	assign X3s2a4 = (~(O5rw84 & Xum2a4));
	assign J3s2a4 = (L4s2a4 & S4s2a4);
	assign S4s2a4 = (~(Yeuw84 & Gwm2a4));
	assign L4s2a4 = (~(M9mw84 & Msm2a4));
	assign Akrx84 = (!Eezx84);
	assign Eezx84 = (~(Z4s2a4 & G5s2a4));
	assign G5s2a4 = (N5s2a4 & U5s2a4);
	assign U5s2a4 = (B6s2a4 & I6s2a4);
	assign I6s2a4 = (P6s2a4 & W6s2a4);
	assign W6s2a4 = (~(I5gw84 & Mlm2a4));
	assign P6s2a4 = (D7s2a4 & K7s2a4);
	assign K7s2a4 = (~(A1yw84 & Hmm2a4));
	assign D7s2a4 = (~(Ckzw84 & Omm2a4));
	assign B6s2a4 = (R7s2a4 & Y7s2a4);
	assign Y7s2a4 = (~(Om9w84 & Jnm2a4));
	assign R7s2a4 = (~(Ashw84 & Qnm2a4));
	assign N5s2a4 = (F8s2a4 & M8s2a4);
	assign M8s2a4 = (T8s2a4 & A9s2a4);
	assign A9s2a4 = (~(G9bw84 & Zom2a4));
	assign T8s2a4 = (~(Yvcw84 & Gpm2a4));
	assign F8s2a4 = (H9s2a4 & O9s2a4);
	assign O9s2a4 = (~(Sejw84 & Bqm2a4));
	assign H9s2a4 = (~(Qiew84 & Iqm2a4));
	assign Z4s2a4 = (V9s2a4 & Cas2a4);
	assign Cas2a4 = (Jas2a4 & Qas2a4);
	assign Qas2a4 = (Xas2a4 & Ebs2a4);
	assign Ebs2a4 = (~(K1lw84 & Fsm2a4));
	assign Xas2a4 = (~(Comw84 & Msm2a4));
	assign Jas2a4 = (Lbs2a4 & Sbs2a4);
	assign Sbs2a4 = (~(Mxpw84 & Htm2a4));
	assign Lbs2a4 = (~(Uaow84 & Otm2a4));
	assign V9s2a4 = (Zbs2a4 & Gcs2a4);
	assign Gcs2a4 = (Ncs2a4 & Ucs2a4);
	assign Ucs2a4 = (~(Ekrw84 & Xum2a4));
	assign Ncs2a4 = (~(W6tw84 & Evm2a4));
	assign Zbs2a4 = (Bds2a4 & Ids2a4);
	assign Ids2a4 = (~(Ggww84 & Zvm2a4));
	assign Bds2a4 = (~(Otuw84 & Gwm2a4));
	assign HWDATA[13] = (!Pds2a4);
	assign Pds2a4 = (Ehm2a4 ? Vw0y84 : Lfrx84);
	assign Vw0y84 = (Wds2a4 & Des2a4);
	assign Des2a4 = (Kes2a4 & Res2a4);
	assign Res2a4 = (Yes2a4 & Ffs2a4);
	assign Ffs2a4 = (~(Xofw84 & Mlm2a4));
	assign Yes2a4 = (Mfs2a4 & Tfs2a4);
	assign Tfs2a4 = (~(Pkxw84 & Hmm2a4));
	assign Mfs2a4 = (~(R3zw84 & Omm2a4));
	assign Kes2a4 = (Ags2a4 & Hgs2a4);
	assign Hgs2a4 = (~(D69w84 & Jnm2a4));
	assign Ags2a4 = (~(Pbhw84 & Qnm2a4));
	assign Wds2a4 = (Ogs2a4 & Vgs2a4);
	assign Vgs2a4 = (Chs2a4 & Jhs2a4);
	assign Jhs2a4 = (~(Hyiw84 & Bqm2a4));
	assign Chs2a4 = (Qhs2a4 & Xhs2a4);
	assign Xhs2a4 = (~(Vsaw84 & Zom2a4));
	assign Qhs2a4 = (~(Nfcw84 & Gpm2a4));
	assign Ogs2a4 = (Dfk2a4 & Eis2a4);
	assign Eis2a4 = (~(F2ew84 & Iqm2a4));
	assign Dfk2a4 = (Lis2a4 & Sis2a4);
	assign Sis2a4 = (Zis2a4 & Gjs2a4);
	assign Gjs2a4 = (Njs2a4 & Ujs2a4);
	assign Ujs2a4 = (~(Zkkw84 & Fsm2a4));
	assign Njs2a4 = (~(R7mw84 & Msm2a4));
	assign Zis2a4 = (Bks2a4 & Iks2a4);
	assign Iks2a4 = (~(Bhpw84 & Htm2a4));
	assign Bks2a4 = (~(Junw84 & Otm2a4));
	assign Lis2a4 = (Pks2a4 & Wks2a4);
	assign Wks2a4 = (Dls2a4 & Kls2a4);
	assign Kls2a4 = (~(T3rw84 & Xum2a4));
	assign Dls2a4 = (~(Lqsw84 & Evm2a4));
	assign Pks2a4 = (Rls2a4 & Yls2a4);
	assign Yls2a4 = (~(Vzvw84 & Zvm2a4));
	assign Rls2a4 = (~(Dduw84 & Gwm2a4));
	assign Lfrx84 = (!Xdzx84);
	assign Xdzx84 = (~(Fms2a4 & Mms2a4));
	assign Mms2a4 = (Tms2a4 & Ans2a4);
	assign Ans2a4 = (Hns2a4 & Ons2a4);
	assign Ons2a4 = (Vns2a4 & Cos2a4);
	assign Cos2a4 = (~(M3gw84 & Mlm2a4));
	assign Vns2a4 = (Jos2a4 & Qos2a4);
	assign Qos2a4 = (~(Ezxw84 & Hmm2a4));
	assign Jos2a4 = (~(Gizw84 & Omm2a4));
	assign Hns2a4 = (Xos2a4 & Eps2a4);
	assign Eps2a4 = (~(Sk9w84 & Jnm2a4));
	assign Xos2a4 = (~(Eqhw84 & Qnm2a4));
	assign Tms2a4 = (Lps2a4 & Sps2a4);
	assign Sps2a4 = (Zps2a4 & Gqs2a4);
	assign Gqs2a4 = (~(K7bw84 & Zom2a4));
	assign Zps2a4 = (~(Cucw84 & Gpm2a4));
	assign Lps2a4 = (Nqs2a4 & Uqs2a4);
	assign Uqs2a4 = (~(Wcjw84 & Bqm2a4));
	assign Nqs2a4 = (~(Ugew84 & Iqm2a4));
	assign Fms2a4 = (Brs2a4 & Irs2a4);
	assign Irs2a4 = (Prs2a4 & Wrs2a4);
	assign Wrs2a4 = (Dss2a4 & Kss2a4);
	assign Kss2a4 = (~(Ozkw84 & Fsm2a4));
	assign Dss2a4 = (~(Gmmw84 & Msm2a4));
	assign Prs2a4 = (Rss2a4 & Yss2a4);
	assign Yss2a4 = (~(Qvpw84 & Htm2a4));
	assign Rss2a4 = (~(Y8ow84 & Otm2a4));
	assign Brs2a4 = (Fts2a4 & Mts2a4);
	assign Mts2a4 = (Tts2a4 & Aus2a4);
	assign Aus2a4 = (~(Iirw84 & Xum2a4));
	assign Tts2a4 = (~(A5tw84 & Evm2a4));
	assign Fts2a4 = (Hus2a4 & Ous2a4);
	assign Ous2a4 = (~(Keww84 & Zvm2a4));
	assign Hus2a4 = (~(Sruw84 & Gwm2a4));
	assign HWDATA[12] = (!Vus2a4);
	assign Vus2a4 = (Ehm2a4 ? W71y84 : B01y84);
	assign W71y84 = (!Shm2a4);
	assign Shm2a4 = (~(Cvs2a4 & Jvs2a4));
	assign Jvs2a4 = (Qvs2a4 & Xvs2a4);
	assign Xvs2a4 = (Ews2a4 & Lws2a4);
	assign Lws2a4 = (~(Cnfw84 & Mlm2a4));
	assign Ews2a4 = (Sws2a4 & Zws2a4);
	assign Zws2a4 = (~(Uixw84 & Hmm2a4));
	assign Sws2a4 = (~(W1zw84 & Omm2a4));
	assign Qvs2a4 = (Gxs2a4 & Nxs2a4);
	assign Nxs2a4 = (~(I49w84 & Jnm2a4));
	assign Gxs2a4 = (~(U9hw84 & Qnm2a4));
	assign Cvs2a4 = (Uxs2a4 & Bys2a4);
	assign Bys2a4 = (Iys2a4 & Pys2a4);
	assign Pys2a4 = (~(Mwiw84 & Bqm2a4));
	assign Iys2a4 = (Wys2a4 & Dzs2a4);
	assign Dzs2a4 = (~(Araw84 & Zom2a4));
	assign Wys2a4 = (~(Sdcw84 & Gpm2a4));
	assign Uxs2a4 = (Sjk2a4 & Kzs2a4);
	assign Kzs2a4 = (~(K0ew84 & Iqm2a4));
	assign Sjk2a4 = (Rzs2a4 & Yzs2a4);
	assign Yzs2a4 = (F0t2a4 & M0t2a4);
	assign M0t2a4 = (T0t2a4 & A1t2a4);
	assign A1t2a4 = (~(Ejkw84 & Fsm2a4));
	assign T0t2a4 = (~(W5mw84 & Msm2a4));
	assign F0t2a4 = (H1t2a4 & O1t2a4);
	assign O1t2a4 = (~(Gfpw84 & Htm2a4));
	assign H1t2a4 = (~(Osnw84 & Otm2a4));
	assign Rzs2a4 = (V1t2a4 & C2t2a4);
	assign C2t2a4 = (J2t2a4 & Q2t2a4);
	assign Q2t2a4 = (~(Y1rw84 & Xum2a4));
	assign J2t2a4 = (~(Qosw84 & Evm2a4));
	assign V1t2a4 = (X2t2a4 & E3t2a4);
	assign E3t2a4 = (~(Ayvw84 & Zvm2a4));
	assign X2t2a4 = (~(Ibuw84 & Gwm2a4));
	assign B01y84 = (L3t2a4 & S3t2a4);
	assign S3t2a4 = (Z3t2a4 & G4t2a4);
	assign G4t2a4 = (N4t2a4 & U4t2a4);
	assign U4t2a4 = (B5t2a4 & I5t2a4);
	assign I5t2a4 = (~(Q1gw84 & Mlm2a4));
	assign B5t2a4 = (P5t2a4 & W5t2a4);
	assign W5t2a4 = (~(Ixxw84 & Hmm2a4));
	assign P5t2a4 = (~(Kgzw84 & Omm2a4));
	assign N4t2a4 = (D6t2a4 & K6t2a4);
	assign K6t2a4 = (~(Wi9w84 & Jnm2a4));
	assign D6t2a4 = (~(Iohw84 & Qnm2a4));
	assign Z3t2a4 = (R6t2a4 & Y6t2a4);
	assign Y6t2a4 = (F7t2a4 & M7t2a4);
	assign M7t2a4 = (~(O5bw84 & Zom2a4));
	assign F7t2a4 = (~(Gscw84 & Gpm2a4));
	assign R6t2a4 = (T7t2a4 & A8t2a4);
	assign A8t2a4 = (~(Abjw84 & Bqm2a4));
	assign T7t2a4 = (~(Yeew84 & Iqm2a4));
	assign L3t2a4 = (H8t2a4 & O8t2a4);
	assign O8t2a4 = (V8t2a4 & C9t2a4);
	assign C9t2a4 = (J9t2a4 & Q9t2a4);
	assign Q9t2a4 = (~(Sxkw84 & Fsm2a4));
	assign J9t2a4 = (~(Kkmw84 & Msm2a4));
	assign V8t2a4 = (X9t2a4 & Eat2a4);
	assign Eat2a4 = (~(Utpw84 & Htm2a4));
	assign X9t2a4 = (~(C7ow84 & Otm2a4));
	assign H8t2a4 = (Lat2a4 & Sat2a4);
	assign Sat2a4 = (Zat2a4 & Gbt2a4);
	assign Gbt2a4 = (~(Mgrw84 & Xum2a4));
	assign Zat2a4 = (~(E3tw84 & Evm2a4));
	assign Lat2a4 = (Nbt2a4 & Ubt2a4);
	assign Ubt2a4 = (~(Ocww84 & Zvm2a4));
	assign Nbt2a4 = (~(Wpuw84 & Gwm2a4));
	assign HWDATA[11] = (Nim2a4 ? Cdzx84 : Yhzx84);
	assign Cdzx84 = (~(Bct2a4 & Ict2a4));
	assign Ict2a4 = (Pct2a4 & Wct2a4);
	assign Wct2a4 = (Ddt2a4 & Kdt2a4);
	assign Kdt2a4 = (Rdt2a4 & Ydt2a4);
	assign Ydt2a4 = (~(Uzfw84 & Mlm2a4));
	assign Rdt2a4 = (Fet2a4 & Met2a4);
	assign Met2a4 = (~(Mvxw84 & Hmm2a4));
	assign Fet2a4 = (~(Oezw84 & Omm2a4));
	assign Ddt2a4 = (Tet2a4 & Aft2a4);
	assign Aft2a4 = (~(Ah9w84 & Jnm2a4));
	assign Tet2a4 = (~(Mmhw84 & Qnm2a4));
	assign Pct2a4 = (Hft2a4 & Oft2a4);
	assign Oft2a4 = (Vft2a4 & Cgt2a4);
	assign Cgt2a4 = (~(S3bw84 & Zom2a4));
	assign Vft2a4 = (~(Kqcw84 & Gpm2a4));
	assign Hft2a4 = (Jgt2a4 & Qgt2a4);
	assign Qgt2a4 = (~(E9jw84 & Bqm2a4));
	assign Jgt2a4 = (~(Cdew84 & Iqm2a4));
	assign Bct2a4 = (Xgt2a4 & Eht2a4);
	assign Eht2a4 = (Lht2a4 & Sht2a4);
	assign Sht2a4 = (Zht2a4 & Git2a4);
	assign Git2a4 = (~(Wvkw84 & Fsm2a4));
	assign Zht2a4 = (~(Oimw84 & Msm2a4));
	assign Lht2a4 = (Nit2a4 & Uit2a4);
	assign Uit2a4 = (~(Yrpw84 & Htm2a4));
	assign Nit2a4 = (~(G5ow84 & Otm2a4));
	assign Xgt2a4 = (Bjt2a4 & Ijt2a4);
	assign Ijt2a4 = (Pjt2a4 & Wjt2a4);
	assign Wjt2a4 = (~(Qerw84 & Xum2a4));
	assign Pjt2a4 = (~(I1tw84 & Evm2a4));
	assign Bjt2a4 = (Dkt2a4 & Kkt2a4);
	assign Kkt2a4 = (~(Saww84 & Zvm2a4));
	assign Dkt2a4 = (~(Aouw84 & Gwm2a4));
	assign Yhzx84 = (~(Rkt2a4 & Ykt2a4));
	assign Ykt2a4 = (Flt2a4 & Mlt2a4);
	assign Mlt2a4 = (Tlt2a4 & Amt2a4);
	assign Amt2a4 = (~(Hlfw84 & Mlm2a4));
	assign Tlt2a4 = (Hmt2a4 & Omt2a4);
	assign Omt2a4 = (~(Zgxw84 & Hmm2a4));
	assign Hmt2a4 = (~(B0zw84 & Omm2a4));
	assign Flt2a4 = (Vmt2a4 & Cnt2a4);
	assign Cnt2a4 = (~(N29w84 & Jnm2a4));
	assign Vmt2a4 = (~(Z7hw84 & Qnm2a4));
	assign Rkt2a4 = (Jnt2a4 & Qnt2a4);
	assign Qnt2a4 = (Xnt2a4 & Eot2a4);
	assign Eot2a4 = (~(Ruiw84 & Bqm2a4));
	assign Xnt2a4 = (Lot2a4 & Sot2a4);
	assign Sot2a4 = (~(Fpaw84 & Zom2a4));
	assign Lot2a4 = (~(Xbcw84 & Gpm2a4));
	assign Jnt2a4 = (~(Hok2a4 | Zot2a4));
	assign Zot2a4 = (Pydw84 & Iqm2a4);
	assign Hok2a4 = (~(Gpt2a4 & Npt2a4));
	assign Npt2a4 = (Upt2a4 & Bqt2a4);
	assign Bqt2a4 = (Iqt2a4 & Pqt2a4);
	assign Pqt2a4 = (~(Jhkw84 & Fsm2a4));
	assign Iqt2a4 = (~(B4mw84 & Msm2a4));
	assign Upt2a4 = (Wqt2a4 & Drt2a4);
	assign Drt2a4 = (~(Ldpw84 & Htm2a4));
	assign Wqt2a4 = (~(Tqnw84 & Otm2a4));
	assign Gpt2a4 = (Krt2a4 & Rrt2a4);
	assign Rrt2a4 = (Yrt2a4 & Fst2a4);
	assign Fst2a4 = (~(D0rw84 & Xum2a4));
	assign Yrt2a4 = (~(Vmsw84 & Evm2a4));
	assign Krt2a4 = (Mst2a4 & Tst2a4);
	assign Tst2a4 = (~(Fwvw84 & Zvm2a4));
	assign Mst2a4 = (~(N9uw84 & Gwm2a4));
	assign HWDATA[10] = (Nim2a4 ? Sezx84 : Rhzx84);
	assign Nim2a4 = (!Ehm2a4);
	assign Ehm2a4 = (Att2a4 & N6r2a4);
	assign Att2a4 = (~(Ralx84 | Htt2a4));
	assign Sezx84 = (~(Ott2a4 & Vtt2a4));
	assign Vtt2a4 = (Cut2a4 & Jut2a4);
	assign Jut2a4 = (Qut2a4 & Xut2a4);
	assign Xut2a4 = (Evt2a4 & Lvt2a4);
	assign Lvt2a4 = (~(Yxfw84 & Mlm2a4));
	assign Evt2a4 = (Svt2a4 & Zvt2a4);
	assign Zvt2a4 = (~(Qtxw84 & Hmm2a4));
	assign Svt2a4 = (~(Sczw84 & Omm2a4));
	assign Qut2a4 = (Gwt2a4 & Nwt2a4);
	assign Nwt2a4 = (~(Ef9w84 & Jnm2a4));
	assign Gwt2a4 = (~(Qkhw84 & Qnm2a4));
	assign Cut2a4 = (Uwt2a4 & Bxt2a4);
	assign Bxt2a4 = (Ixt2a4 & Pxt2a4);
	assign Pxt2a4 = (~(W1bw84 & Zom2a4));
	assign Ixt2a4 = (~(Oocw84 & Gpm2a4));
	assign Uwt2a4 = (Wxt2a4 & Dyt2a4);
	assign Dyt2a4 = (~(I7jw84 & Bqm2a4));
	assign Wxt2a4 = (~(Gbew84 & Iqm2a4));
	assign Ott2a4 = (Kyt2a4 & Ryt2a4);
	assign Ryt2a4 = (Yyt2a4 & Fzt2a4);
	assign Fzt2a4 = (Mzt2a4 & Tzt2a4);
	assign Tzt2a4 = (~(Aukw84 & Fsm2a4));
	assign Mzt2a4 = (~(Sgmw84 & Msm2a4));
	assign Yyt2a4 = (A0u2a4 & H0u2a4);
	assign H0u2a4 = (~(Cqpw84 & Htm2a4));
	assign A0u2a4 = (~(K3ow84 & Otm2a4));
	assign Kyt2a4 = (O0u2a4 & V0u2a4);
	assign V0u2a4 = (C1u2a4 & J1u2a4);
	assign J1u2a4 = (~(Ucrw84 & Xum2a4));
	assign C1u2a4 = (~(Mzsw84 & Evm2a4));
	assign O0u2a4 = (Q1u2a4 & X1u2a4);
	assign X1u2a4 = (~(W8ww84 & Zvm2a4));
	assign Q1u2a4 = (~(Emuw84 & Gwm2a4));
	assign Rhzx84 = (~(E2u2a4 & L2u2a4));
	assign L2u2a4 = (S2u2a4 & Z2u2a4);
	assign Z2u2a4 = (G3u2a4 & N3u2a4);
	assign N3u2a4 = (~(Mjfw84 & Mlm2a4));
	assign G3u2a4 = (U3u2a4 & B4u2a4);
	assign B4u2a4 = (~(Efxw84 & Hmm2a4));
	assign Hmm2a4 = (I4u2a4 & Mdxw84);
	assign I4u2a4 = (~(P4u2a4 | W4u2a4));
	assign U3u2a4 = (~(Gyyw84 & Omm2a4));
	assign Omm2a4 = (D5u2a4 & K5u2a4);
	assign D5u2a4 = (~(W4u2a4 | Mdxw84));
	assign S2u2a4 = (R5u2a4 & Y5u2a4);
	assign Y5u2a4 = (~(S09w84 & Jnm2a4));
	assign R5u2a4 = (~(E6hw84 & Qnm2a4));
	assign E2u2a4 = (F6u2a4 & M6u2a4);
	assign M6u2a4 = (T6u2a4 & A7u2a4);
	assign A7u2a4 = (~(Wsiw84 & Bqm2a4));
	assign T6u2a4 = (H7u2a4 & O7u2a4);
	assign O7u2a4 = (~(Knaw84 & Zom2a4));
	assign H7u2a4 = (~(Cacw84 & Gpm2a4));
	assign F6u2a4 = (Mnk2a4 & V7u2a4);
	assign V7u2a4 = (~(Uwdw84 & Iqm2a4));
	assign Mnk2a4 = (C8u2a4 & J8u2a4);
	assign J8u2a4 = (Q8u2a4 & X8u2a4);
	assign X8u2a4 = (E9u2a4 & L9u2a4);
	assign L9u2a4 = (~(Ofkw84 & Fsm2a4));
	assign E9u2a4 = (~(G2mw84 & Msm2a4));
	assign Q8u2a4 = (S9u2a4 & Z9u2a4);
	assign Z9u2a4 = (~(Qbpw84 & Htm2a4));
	assign S9u2a4 = (~(Yonw84 & Otm2a4));
	assign C8u2a4 = (Gau2a4 & Nau2a4);
	assign Nau2a4 = (Uau2a4 & Bbu2a4);
	assign Bbu2a4 = (~(Iyqw84 & Xum2a4));
	assign Uau2a4 = (~(Alsw84 & Evm2a4));
	assign Gau2a4 = (Ibu2a4 & Pbu2a4);
	assign Pbu2a4 = (~(Kuvw84 & Zvm2a4));
	assign Ibu2a4 = (~(S7uw84 & Gwm2a4));
	assign HWDATA[0] = (~(Ralx84 | Yn0y84));
	assign Yn0y84 = (!Vghx84);
	assign Vghx84 = (~(Wbu2a4 & Dcu2a4));
	assign Dcu2a4 = (Kcu2a4 & Rcu2a4);
	assign Rcu2a4 = (Ycu2a4 & Fdu2a4);
	assign Fdu2a4 = (~(Wffw84 & Mlm2a4));
	assign Mlm2a4 = (~(Mdu2a4 | Tdu2a4));
	assign Ycu2a4 = (~(Cx8w84 & Jnm2a4));
	assign Jnm2a4 = (~(Aeu2a4 | W4u2a4));
	assign Kcu2a4 = (Heu2a4 & Oeu2a4);
	assign Oeu2a4 = (~(O2hw84 & Qnm2a4));
	assign Qnm2a4 = (~(Mdu2a4 | P4u2a4));
	assign Heu2a4 = (~(Ujaw84 & Zom2a4));
	assign Zom2a4 = (~(Tdu2a4 | W4u2a4));
	assign Wbu2a4 = (Veu2a4 & Cfu2a4);
	assign Cfu2a4 = (Jfu2a4 & Qfu2a4);
	assign Qfu2a4 = (~(M6cw84 & Gpm2a4));
	assign Gpm2a4 = (~(Xfu2a4 | W4u2a4));
	assign W4u2a4 = (S4vx84 | Zxux84);
	assign Jfu2a4 = (~(Gpiw84 & Bqm2a4));
	assign Bqm2a4 = (~(Xfu2a4 | Mdu2a4));
	assign Veu2a4 = (Wlk2a4 & Egu2a4);
	assign Egu2a4 = (~(Etdw84 & Iqm2a4));
	assign Iqm2a4 = (~(Aeu2a4 | Mdu2a4));
	assign Mdu2a4 = (S4vx84 | Ab5w84);
	assign S4vx84 = (!Tc5w84);
	assign Wlk2a4 = (Lgu2a4 & Sgu2a4);
	assign Sgu2a4 = (Zgu2a4 & Ghu2a4);
	assign Ghu2a4 = (Nhu2a4 & Uhu2a4);
	assign Uhu2a4 = (~(Ybkw84 & Fsm2a4));
	assign Fsm2a4 = (~(Biu2a4 | Aeu2a4));
	assign Nhu2a4 = (~(Qylw84 & Msm2a4));
	assign Msm2a4 = (~(Biu2a4 | Tdu2a4));
	assign Zgu2a4 = (Iiu2a4 & Piu2a4);
	assign Piu2a4 = (~(A8pw84 & Htm2a4));
	assign Htm2a4 = (~(Biu2a4 | Xfu2a4));
	assign Iiu2a4 = (~(Ilnw84 & Otm2a4));
	assign Otm2a4 = (~(Biu2a4 | P4u2a4));
	assign Biu2a4 = (Zxux84 | Tc5w84);
	assign Zxux84 = (!Ab5w84);
	assign Lgu2a4 = (Wiu2a4 & Dju2a4);
	assign Dju2a4 = (Kju2a4 & Rju2a4);
	assign Rju2a4 = (~(Suqw84 & Xum2a4));
	assign Xum2a4 = (~(Yju2a4 | Aeu2a4));
	assign Aeu2a4 = (Oghx84 | Q3vx84);
	assign Kju2a4 = (~(Khsw84 & Evm2a4));
	assign Evm2a4 = (~(Yju2a4 | Tdu2a4));
	assign Tdu2a4 = (Oghx84 | O75w84);
	assign Oghx84 = (!H95w84);
	assign Wiu2a4 = (Fku2a4 & Mku2a4);
	assign Mku2a4 = (~(Uqvw84 & Zvm2a4));
	assign Zvm2a4 = (~(Yju2a4 | Xfu2a4));
	assign Xfu2a4 = (O75w84 | H95w84);
	assign Fku2a4 = (~(C4uw84 & Gwm2a4));
	assign Gwm2a4 = (~(Yju2a4 | P4u2a4));
	assign P4u2a4 = (!K5u2a4);
	assign K5u2a4 = (~(Q3vx84 | H95w84));
	assign Q3vx84 = (!O75w84);
	assign Yju2a4 = (Ab5w84 | Tc5w84);
	assign Ralx84 = (!C45w84);
	assign HTRANS[1] = (Nna2a4 ? HPROT[3] : Tku2a4);
	assign Nna2a4 = (~(Alu2a4 | HPROT[0]));
	assign Tku2a4 = (Hlu2a4 & Olu2a4);
	assign Olu2a4 = (Vlu2a4 & Dkix84);
	assign Vlu2a4 = (~(M1hx84 | Y0hx84));
	assign M1hx84 = (Cmu2a4 & Jmu2a4);
	assign Jmu2a4 = (~(Cza2a4 & Qmu2a4));
	assign Qmu2a4 = (Xmu2a4 | Nqvx84);
	assign Nqvx84 = (!Oya2a4);
	assign Cmu2a4 = (~(Xmu2a4 & N1p2a4));
	assign Hlu2a4 = (O2hx84 & Enu2a4);
	assign Enu2a4 = (A2hx84 | HADDR[28]);
	assign A2hx84 = (~(Lnu2a4 & HADDR[29]));
	assign Lnu2a4 = (HADDR[31] & HADDR[30]);
	assign HSIZE[1] = (~(Alu2a4 & Snu2a4));
	assign Snu2a4 = (F1hx84 | N6r2a4);
	assign HSIZE[0] = (Znu2a4 & Htt2a4);
	assign Znu2a4 = (Alu2a4 & Dkix84);
	assign HPROT[3] = (~(HPROT[2] & Gou2a4));
	assign Gou2a4 = (Nou2a4 | HADDR[31]);
	assign Nou2a4 = (!HADDR[29]);
	assign HPROT[2] = (HADDR[29] | HADDR[30]);
	assign HPROT[0] = (~(Uou2a4 & Bpu2a4));
	assign Bpu2a4 = (Ipu2a4 & Ppu2a4);
	assign Ppu2a4 = (Wpu2a4 & Fem2a4);
	assign Fem2a4 = (~(Dqu2a4 & Krix84));
	assign Dqu2a4 = (~(Mycx84 | D53x84));
	assign Mycx84 = (!M0px84);
	assign Wpu2a4 = (~(Kqu2a4 & Rqu2a4));
	assign Rqu2a4 = (~(Xcmx84 | Wqbx84));
	assign Kqu2a4 = (Laix84 & F2gx84);
	assign Ipu2a4 = (Yqu2a4 & Fru2a4);
	assign Fru2a4 = (~(Mru2a4 & U8lx84));
	assign U8lx84 = (Pz2x84 & Qxmx84);
	assign Mru2a4 = (~(N4bx84 | Ambx84));
	assign Yqu2a4 = (~(Tru2a4 & Hgvx84));
	assign Tru2a4 = (~(Asu2a4 & Hsu2a4));
	assign Hsu2a4 = (~(Osu2a4 & Qxmx84));
	assign Osu2a4 = (~(Vsu2a4 & Ctu2a4));
	assign Ctu2a4 = (N4bx84 | Rybx84);
	assign Vsu2a4 = (S1dx84 | Pz2x84);
	assign Asu2a4 = (Nbix84 | N052a4);
	assign Uou2a4 = (Jtu2a4 & Qtu2a4);
	assign Qtu2a4 = (Xtu2a4 & Euu2a4);
	assign Euu2a4 = (~(Luu2a4 & H6dx84));
	assign Luu2a4 = (~(Mf72a4 & Suu2a4));
	assign Suu2a4 = (~(Zuu2a4 & Phdx84));
	assign Zuu2a4 = (Laix84 & Drbx84);
	assign Mf72a4 = (A1px84 & Gvu2a4);
	assign Gvu2a4 = (~(Nvu2a4 & Rzhx84));
	assign Nvu2a4 = (Uacx84 & G4bx84);
	assign A1px84 = (Vfwx84 | Ucox84);
	assign Vfwx84 = (!Aq42a4);
	assign Xtu2a4 = (~(Fo52a4 & Mlbx84));
	assign Fo52a4 = (Lw72a4 & Pz2x84);
	assign Jtu2a4 = (Uvu2a4 & Bwu2a4);
	assign Bwu2a4 = (~(Uacx84 & A7cx84));
	assign HADDR[9] = (~(Iwu2a4 & Pwu2a4));
	assign Pwu2a4 = (~(Ao63a4[8] & F1hx84));
	assign Iwu2a4 = (Wwu2a4 & Dxu2a4);
	assign Dxu2a4 = (Kxu2a4 | Rsax84);
	assign Rsax84 = (!Xb1y84);
	assign Xb1y84 = (~(Rxu2a4 & Yxu2a4));
	assign Yxu2a4 = (~(Ob9w84 & M7ix84));
	assign Rxu2a4 = (Fyu2a4 & Myu2a4);
	assign Myu2a4 = (~(Tyu2a4 & Azu2a4));
	assign Azu2a4 = (~(Hzu2a4 & Ozu2a4));
	assign Ozu2a4 = (Vzu2a4 & C0v2a4);
	assign C0v2a4 = (J0v2a4 & Q0v2a4);
	assign Q0v2a4 = (~(Tmcw84 & X0v2a4));
	assign J0v2a4 = (E1v2a4 & L1v2a4);
	assign L1v2a4 = (~(Vrxw84 & S1v2a4));
	assign E1v2a4 = (~(Xazw84 & Z1v2a4));
	assign Vzu2a4 = (G2v2a4 & N2v2a4);
	assign N2v2a4 = (~(Dwfw84 & U2v2a4));
	assign G2v2a4 = (~(L9ew84 & B3v2a4));
	assign Hzu2a4 = (I3v2a4 & P3v2a4);
	assign P3v2a4 = (W3v2a4 & D4v2a4);
	assign D4v2a4 = (~(N5jw84 & K4v2a4));
	assign W3v2a4 = (~(Vihw84 & R4v2a4));
	assign I3v2a4 = (~(Fdg2a4 | Y4v2a4));
	assign Y4v2a4 = (B0bw84 & F5v2a4);
	assign Fyu2a4 = (~(Jd9w84 & M5v2a4));
	assign Wwu2a4 = (~(T5v2a4 & Qp63a4[9]));
	assign HADDR[8] = (~(A6v2a4 & H6v2a4));
	assign H6v2a4 = (~(Ao63a4[7] & F1hx84));
	assign A6v2a4 = (O6v2a4 & V6v2a4);
	assign V6v2a4 = (Kxu2a4 | Ysax84);
	assign Ysax84 = (!H31y84);
	assign H31y84 = (~(C7v2a4 & J7v2a4));
	assign J7v2a4 = (~(T99w84 & M7ix84));
	assign C7v2a4 = (Q7v2a4 & X7v2a4);
	assign X7v2a4 = (~(Tyu2a4 & E8v2a4));
	assign E8v2a4 = (~(L8v2a4 & S8v2a4));
	assign S8v2a4 = (Z8v2a4 & G9v2a4);
	assign G9v2a4 = (N9v2a4 & U9v2a4);
	assign U9v2a4 = (~(Ykcw84 & X0v2a4));
	assign N9v2a4 = (Bav2a4 & Iav2a4);
	assign Iav2a4 = (~(Aqxw84 & S1v2a4));
	assign Bav2a4 = (~(C9zw84 & Z1v2a4));
	assign Z8v2a4 = (Pav2a4 & Wav2a4);
	assign Wav2a4 = (~(Iufw84 & U2v2a4));
	assign Pav2a4 = (~(Q7ew84 & B3v2a4));
	assign L8v2a4 = (Dbv2a4 & Kbv2a4);
	assign Kbv2a4 = (Rbv2a4 & Ybv2a4);
	assign Ybv2a4 = (~(S3jw84 & K4v2a4));
	assign Rbv2a4 = (~(Ahhw84 & R4v2a4));
	assign Dbv2a4 = (~(Bxf2a4 | Fcv2a4));
	assign Fcv2a4 = (Gyaw84 & F5v2a4);
	assign Q7v2a4 = (~(Ob9w84 & M5v2a4));
	assign O6v2a4 = (~(T5v2a4 & Qp63a4[8]));
	assign HADDR[7] = (~(Mcv2a4 & Tcv2a4));
	assign Tcv2a4 = (~(Ao63a4[6] & F1hx84));
	assign Mcv2a4 = (Adv2a4 & Hdv2a4);
	assign Hdv2a4 = (Kxu2a4 | Ftax84);
	assign Ftax84 = (!Dazx84);
	assign Dazx84 = (~(Odv2a4 & Vdv2a4));
	assign Vdv2a4 = (~(Y79w84 & M7ix84));
	assign Odv2a4 = (Cev2a4 & Jev2a4);
	assign Jev2a4 = (~(Tyu2a4 & Qev2a4));
	assign Qev2a4 = (~(Xev2a4 & Efv2a4));
	assign Efv2a4 = (Lfv2a4 & Sfv2a4);
	assign Sfv2a4 = (Zfv2a4 & Ggv2a4);
	assign Ggv2a4 = (~(X0v2a4 & Djcw84));
	assign Zfv2a4 = (Ngv2a4 & Ugv2a4);
	assign Ugv2a4 = (~(S1v2a4 & Foxw84));
	assign Ngv2a4 = (~(Z1v2a4 & H7zw84));
	assign Lfv2a4 = (Bhv2a4 & Ihv2a4);
	assign Ihv2a4 = (~(U2v2a4 & Nsfw84));
	assign Bhv2a4 = (~(B3v2a4 & V5ew84));
	assign Xev2a4 = (Phv2a4 & Whv2a4);
	assign Whv2a4 = (Div2a4 & Kiv2a4);
	assign Kiv2a4 = (~(K4v2a4 & X1jw84));
	assign Div2a4 = (~(R4v2a4 & Ffhw84));
	assign Phv2a4 = (~(Dyf2a4 | Riv2a4));
	assign Riv2a4 = (F5v2a4 & Lwaw84);
	assign Cev2a4 = (~(M5v2a4 & T99w84));
	assign Adv2a4 = (~(Qp63a4[7] & T5v2a4));
	assign HADDR[6] = (~(Yiv2a4 & Fjv2a4));
	assign Fjv2a4 = (~(Ao63a4[5] & F1hx84));
	assign Yiv2a4 = (Mjv2a4 & Tjv2a4);
	assign Tjv2a4 = (Kxu2a4 | Mtax84);
	assign Mtax84 = (Akv2a4 & Hkv2a4);
	assign Hkv2a4 = (~(D69w84 & M7ix84));
	assign Akv2a4 = (Okv2a4 & Vkv2a4);
	assign Vkv2a4 = (~(Tyu2a4 & Clv2a4));
	assign Clv2a4 = (~(Jlv2a4 & Qlv2a4));
	assign Qlv2a4 = (Xlv2a4 & Emv2a4);
	assign Emv2a4 = (Lmv2a4 & Smv2a4);
	assign Smv2a4 = (~(Ihcw84 & X0v2a4));
	assign Lmv2a4 = (Zmv2a4 & Gnv2a4);
	assign Gnv2a4 = (~(Kmxw84 & S1v2a4));
	assign Zmv2a4 = (~(M5zw84 & Z1v2a4));
	assign Xlv2a4 = (Nnv2a4 & Unv2a4);
	assign Unv2a4 = (~(Sqfw84 & U2v2a4));
	assign Nnv2a4 = (~(A4ew84 & B3v2a4));
	assign Jlv2a4 = (Bov2a4 & Iov2a4);
	assign Iov2a4 = (Pov2a4 & Wov2a4);
	assign Wov2a4 = (~(C0jw84 & K4v2a4));
	assign Pov2a4 = (~(Kdhw84 & R4v2a4));
	assign Bov2a4 = (~(Ixf2a4 | Dpv2a4));
	assign Dpv2a4 = (Quaw84 & F5v2a4);
	assign Okv2a4 = (~(Y79w84 & M5v2a4));
	assign Mjv2a4 = (~(T5v2a4 & Qp63a4[6]));
	assign HADDR[5] = (~(Kpv2a4 & Rpv2a4));
	assign Rpv2a4 = (~(Ao63a4[4] & F1hx84));
	assign Kpv2a4 = (Ypv2a4 & Fqv2a4);
	assign Fqv2a4 = (Kxu2a4 | Ttax84);
	assign Ttax84 = (!Ly0y84);
	assign Ly0y84 = (~(Mqv2a4 & Tqv2a4));
	assign Tqv2a4 = (~(I49w84 & M7ix84));
	assign Mqv2a4 = (Arv2a4 & Hrv2a4);
	assign Hrv2a4 = (~(Tyu2a4 & Orv2a4));
	assign Orv2a4 = (~(Vrv2a4 & Csv2a4));
	assign Csv2a4 = (Jsv2a4 & Qsv2a4);
	assign Qsv2a4 = (Xsv2a4 & Etv2a4);
	assign Etv2a4 = (~(Nfcw84 & X0v2a4));
	assign Xsv2a4 = (Ltv2a4 & Stv2a4);
	assign Stv2a4 = (~(Pkxw84 & S1v2a4));
	assign Ltv2a4 = (~(R3zw84 & Z1v2a4));
	assign Jsv2a4 = (Ztv2a4 & Guv2a4);
	assign Guv2a4 = (~(Xofw84 & U2v2a4));
	assign Ztv2a4 = (~(F2ew84 & B3v2a4));
	assign Vrv2a4 = (Nuv2a4 & Uuv2a4);
	assign Uuv2a4 = (Bvv2a4 & Ivv2a4);
	assign Ivv2a4 = (~(Hyiw84 & K4v2a4));
	assign Bvv2a4 = (~(Pbhw84 & R4v2a4));
	assign Nuv2a4 = (~(Kyf2a4 | Pvv2a4));
	assign Pvv2a4 = (Vsaw84 & F5v2a4);
	assign Arv2a4 = (~(D69w84 & M5v2a4));
	assign Ypv2a4 = (~(T5v2a4 & Qp63a4[5]));
	assign HADDR[4] = (~(Wvv2a4 & Dwv2a4));
	assign Dwv2a4 = (~(Ao63a4[3] & F1hx84));
	assign Wvv2a4 = (Kwv2a4 & Rwv2a4);
	assign Rwv2a4 = (Kxu2a4 | Auax84);
	assign Auax84 = (!M91y84);
	assign M91y84 = (~(Ywv2a4 & Fxv2a4));
	assign Fxv2a4 = (~(N29w84 & M7ix84));
	assign Ywv2a4 = (Mxv2a4 & Txv2a4);
	assign Txv2a4 = (~(Tyu2a4 & Ayv2a4));
	assign Ayv2a4 = (~(Hyv2a4 & Oyv2a4));
	assign Oyv2a4 = (Vyv2a4 & Czv2a4);
	assign Czv2a4 = (Jzv2a4 & Qzv2a4);
	assign Qzv2a4 = (~(Sdcw84 & X0v2a4));
	assign Jzv2a4 = (Xzv2a4 & E0w2a4);
	assign E0w2a4 = (~(Uixw84 & S1v2a4));
	assign Xzv2a4 = (~(W1zw84 & Z1v2a4));
	assign Vyv2a4 = (L0w2a4 & S0w2a4);
	assign S0w2a4 = (~(Cnfw84 & U2v2a4));
	assign L0w2a4 = (~(K0ew84 & B3v2a4));
	assign Hyv2a4 = (Z0w2a4 & G1w2a4);
	assign G1w2a4 = (N1w2a4 & U1w2a4);
	assign U1w2a4 = (~(Mwiw84 & K4v2a4));
	assign N1w2a4 = (~(U9hw84 & R4v2a4));
	assign Z0w2a4 = (~(Otf2a4 | B2w2a4));
	assign B2w2a4 = (Araw84 & F5v2a4);
	assign Mxv2a4 = (~(I49w84 & M5v2a4));
	assign Kwv2a4 = (~(T5v2a4 & Qp63a4[4]));
	assign HADDR[3] = (~(I2w2a4 & P2w2a4));
	assign P2w2a4 = (~(Ao63a4[2] & F1hx84));
	assign I2w2a4 = (W2w2a4 & D3w2a4);
	assign D3w2a4 = (Kxu2a4 | Huax84);
	assign Huax84 = (!Bm0y84);
	assign Bm0y84 = (~(K3w2a4 & R3w2a4));
	assign R3w2a4 = (~(S09w84 & M7ix84));
	assign K3w2a4 = (Y3w2a4 & F4w2a4);
	assign F4w2a4 = (~(Tyu2a4 & M4w2a4));
	assign M4w2a4 = (~(T4w2a4 & A5w2a4));
	assign A5w2a4 = (H5w2a4 & O5w2a4);
	assign O5w2a4 = (V5w2a4 & C6w2a4);
	assign C6w2a4 = (~(Xbcw84 & X0v2a4));
	assign V5w2a4 = (J6w2a4 & Q6w2a4);
	assign Q6w2a4 = (~(Zgxw84 & S1v2a4));
	assign J6w2a4 = (~(B0zw84 & Z1v2a4));
	assign H5w2a4 = (X6w2a4 & E7w2a4);
	assign E7w2a4 = (~(Hlfw84 & U2v2a4));
	assign X6w2a4 = (~(Pydw84 & B3v2a4));
	assign T4w2a4 = (L7w2a4 & S7w2a4);
	assign S7w2a4 = (Z7w2a4 & G8w2a4);
	assign G8w2a4 = (~(Ruiw84 & K4v2a4));
	assign Z7w2a4 = (~(Z7hw84 & R4v2a4));
	assign L7w2a4 = (~(Xuf2a4 | N8w2a4));
	assign N8w2a4 = (Fpaw84 & F5v2a4);
	assign Y3w2a4 = (~(N29w84 & M5v2a4));
	assign W2w2a4 = (~(Qp63a4[3] & T5v2a4));
	assign HADDR[31] = (~(U8w2a4 & B9w2a4));
	assign B9w2a4 = (~(Ao63a4[30] & F1hx84));
	assign U8w2a4 = (I9w2a4 & P9w2a4);
	assign P9w2a4 = (Kxu2a4 | J32y84);
	assign J32y84 = (!O7xx84);
	assign O7xx84 = (~(W9w2a4 & Daw2a4));
	assign Daw2a4 = (~(Cgaw84 & M7ix84));
	assign W9w2a4 = (Kaw2a4 & Raw2a4);
	assign Raw2a4 = (~(Tyu2a4 & Yaw2a4));
	assign Yaw2a4 = (~(Fbw2a4 & Mbw2a4));
	assign Mbw2a4 = (Tbw2a4 & Acw2a4);
	assign Acw2a4 = (Hcw2a4 & Ocw2a4);
	assign Ocw2a4 = (~(X0v2a4 & Irdw84));
	assign Hcw2a4 = (Vcw2a4 & Cdw2a4);
	assign Cdw2a4 = (~(S1v2a4 & Kwyw84));
	assign Vcw2a4 = (~(Z1v2a4 & Mf0x84));
	assign Tbw2a4 = (Jdw2a4 & Qdw2a4);
	assign Qdw2a4 = (~(U2v2a4 & S0hw84));
	assign Jdw2a4 = (~(B3v2a4 & Aefw84));
	assign Fbw2a4 = (Xdw2a4 & Eew2a4);
	assign Eew2a4 = (Lew2a4 & Sew2a4);
	assign Sew2a4 = (~(K4v2a4 & Cakw84));
	assign Lew2a4 = (~(R4v2a4 & Kniw84));
	assign Xdw2a4 = (~(K5g2a4 | Zew2a4));
	assign Zew2a4 = (F5v2a4 & Q4cw84);
	assign Kaw2a4 = (~(M5v2a4 & Yhaw84));
	assign I9w2a4 = (~(T5v2a4 & Qp63a4[31]));
	assign HADDR[30] = (~(Gfw2a4 & Nfw2a4));
	assign Nfw2a4 = (~(Ao63a4[29] & F1hx84));
	assign Gfw2a4 = (Ufw2a4 & Bgw2a4);
	assign Bgw2a4 = (Kxu2a4 | Ouax84);
	assign Ouax84 = (!Zj1y84);
	assign Zj1y84 = (~(Igw2a4 & Pgw2a4));
	assign Pgw2a4 = (~(Geaw84 & M7ix84));
	assign Igw2a4 = (Wgw2a4 & Dhw2a4);
	assign Dhw2a4 = (~(Tyu2a4 & Khw2a4));
	assign Khw2a4 = (~(Rhw2a4 & Yhw2a4));
	assign Yhw2a4 = (Fiw2a4 & Miw2a4);
	assign Miw2a4 = (Tiw2a4 & Ajw2a4);
	assign Ajw2a4 = (~(Mpdw84 & X0v2a4));
	assign Tiw2a4 = (Hjw2a4 & Ojw2a4);
	assign Ojw2a4 = (~(Ouyw84 & S1v2a4));
	assign Hjw2a4 = (~(Qd0x84 & Z1v2a4));
	assign Fiw2a4 = (Vjw2a4 & Ckw2a4);
	assign Ckw2a4 = (~(Wygw84 & U2v2a4));
	assign Vjw2a4 = (~(Ecfw84 & B3v2a4));
	assign Rhw2a4 = (Jkw2a4 & Qkw2a4);
	assign Qkw2a4 = (Xkw2a4 & Elw2a4);
	assign Elw2a4 = (~(G8kw84 & K4v2a4));
	assign Xkw2a4 = (~(Oliw84 & R4v2a4));
	assign Jkw2a4 = (~(P4g2a4 | Llw2a4));
	assign Llw2a4 = (U2cw84 & F5v2a4);
	assign Wgw2a4 = (~(Cgaw84 & M5v2a4));
	assign Ufw2a4 = (~(T5v2a4 & Qp63a4[30]));
	assign HADDR[2] = (~(Slw2a4 & Zlw2a4));
	assign Zlw2a4 = (~(Qp63a4[2] & T5v2a4));
	assign Slw2a4 = (Gmw2a4 & Nmw2a4);
	assign Nmw2a4 = (~(F1hx84 & Umw2a4));
	assign Umw2a4 = (Bnw2a4 ^ Wrax84);
	assign Wrax84 = (Dsax84 ^ V55w84);
	assign Bnw2a4 = (Tk63a4[0] & Prax84);
	assign Gmw2a4 = (Kxu2a4 | Lwax84);
	assign Lwax84 = (!Ascx84);
	assign Ascx84 = (~(Inw2a4 & Pnw2a4));
	assign Pnw2a4 = (~(Xy8w84 & M7ix84));
	assign Inw2a4 = (Wnw2a4 & Dow2a4);
	assign Dow2a4 = (~(Tyu2a4 & Kow2a4));
	assign Kow2a4 = (~(Row2a4 & Yow2a4));
	assign Yow2a4 = (Fpw2a4 & Mpw2a4);
	assign Mpw2a4 = (Tpw2a4 & Aqw2a4);
	assign Aqw2a4 = (~(Cacw84 & X0v2a4));
	assign Tpw2a4 = (Hqw2a4 & Oqw2a4);
	assign Oqw2a4 = (~(Efxw84 & S1v2a4));
	assign Hqw2a4 = (~(Gyyw84 & Z1v2a4));
	assign Fpw2a4 = (Vqw2a4 & Crw2a4);
	assign Crw2a4 = (~(Mjfw84 & U2v2a4));
	assign Vqw2a4 = (~(Uwdw84 & B3v2a4));
	assign Row2a4 = (Jrw2a4 & Qrw2a4);
	assign Qrw2a4 = (Xrw2a4 & Esw2a4);
	assign Esw2a4 = (~(Wsiw84 & K4v2a4));
	assign Xrw2a4 = (~(E6hw84 & R4v2a4));
	assign Jrw2a4 = (~(Vtf2a4 | Lsw2a4));
	assign Lsw2a4 = (Knaw84 & F5v2a4);
	assign Wnw2a4 = (~(S09w84 & M5v2a4));
	assign HADDR[29] = (~(Ssw2a4 & Zsw2a4));
	assign Zsw2a4 = (~(Ao63a4[28] & F1hx84));
	assign Ssw2a4 = (Gtw2a4 & Ntw2a4);
	assign Ntw2a4 = (Kxu2a4 | Swax84);
	assign Swax84 = (!Rm1y84);
	assign Rm1y84 = (~(Utw2a4 & Buw2a4));
	assign Buw2a4 = (~(Kcaw84 & M7ix84));
	assign Utw2a4 = (Iuw2a4 & Puw2a4);
	assign Puw2a4 = (~(Tyu2a4 & Wuw2a4));
	assign Wuw2a4 = (~(Dvw2a4 & Kvw2a4));
	assign Kvw2a4 = (Rvw2a4 & Yvw2a4);
	assign Yvw2a4 = (Fww2a4 & Mww2a4);
	assign Mww2a4 = (~(Qndw84 & X0v2a4));
	assign Fww2a4 = (Tww2a4 & Axw2a4);
	assign Axw2a4 = (~(Ssyw84 & S1v2a4));
	assign Tww2a4 = (~(Ub0x84 & Z1v2a4));
	assign Rvw2a4 = (Hxw2a4 & Oxw2a4);
	assign Oxw2a4 = (~(Axgw84 & U2v2a4));
	assign Hxw2a4 = (~(Iafw84 & B3v2a4));
	assign Dvw2a4 = (Vxw2a4 & Cyw2a4);
	assign Cyw2a4 = (Jyw2a4 & Qyw2a4);
	assign Qyw2a4 = (~(K6kw84 & K4v2a4));
	assign Jyw2a4 = (~(Sjiw84 & R4v2a4));
	assign Vxw2a4 = (~(R5g2a4 | Xyw2a4));
	assign Xyw2a4 = (Y0cw84 & F5v2a4);
	assign Iuw2a4 = (~(Geaw84 & M5v2a4));
	assign Gtw2a4 = (~(T5v2a4 & Qp63a4[29]));
	assign HADDR[28] = (~(Ezw2a4 & Lzw2a4));
	assign Lzw2a4 = (~(Ao63a4[27] & F1hx84));
	assign Ezw2a4 = (Szw2a4 & Zzw2a4);
	assign Zzw2a4 = (Kxu2a4 | Zwax84);
	assign Zwax84 = (!R90y84);
	assign R90y84 = (~(G0x2a4 & N0x2a4));
	assign N0x2a4 = (~(Oaaw84 & M7ix84));
	assign G0x2a4 = (U0x2a4 & B1x2a4);
	assign B1x2a4 = (~(Tyu2a4 & I1x2a4));
	assign I1x2a4 = (~(P1x2a4 & W1x2a4));
	assign W1x2a4 = (D2x2a4 & K2x2a4);
	assign K2x2a4 = (R2x2a4 & Y2x2a4);
	assign Y2x2a4 = (~(Uldw84 & X0v2a4));
	assign R2x2a4 = (F3x2a4 & M3x2a4);
	assign M3x2a4 = (~(Wqyw84 & S1v2a4));
	assign F3x2a4 = (~(Y90x84 & Z1v2a4));
	assign D2x2a4 = (T3x2a4 & A4x2a4);
	assign A4x2a4 = (~(Evgw84 & U2v2a4));
	assign T3x2a4 = (~(M8fw84 & B3v2a4));
	assign P1x2a4 = (H4x2a4 & O4x2a4);
	assign O4x2a4 = (V4x2a4 & C5x2a4);
	assign C5x2a4 = (~(O4kw84 & K4v2a4));
	assign V4x2a4 = (~(Whiw84 & R4v2a4));
	assign H4x2a4 = (~(A7g2a4 | J5x2a4));
	assign J5x2a4 = (Czbw84 & F5v2a4);
	assign U0x2a4 = (~(Kcaw84 & M5v2a4));
	assign Szw2a4 = (~(Qp63a4[28] & T5v2a4));
	assign HADDR[27] = (~(Q5x2a4 & X5x2a4));
	assign X5x2a4 = (~(Ao63a4[26] & F1hx84));
	assign Q5x2a4 = (E6x2a4 & L6x2a4);
	assign L6x2a4 = (Kxu2a4 | Gxax84);
	assign Gxax84 = (!Jzyx84);
	assign Jzyx84 = (~(S6x2a4 & Z6x2a4));
	assign Z6x2a4 = (~(S8aw84 & M7ix84));
	assign S6x2a4 = (G7x2a4 & N7x2a4);
	assign N7x2a4 = (~(Tyu2a4 & U7x2a4));
	assign U7x2a4 = (~(B8x2a4 & I8x2a4));
	assign I8x2a4 = (P8x2a4 & W8x2a4);
	assign W8x2a4 = (D9x2a4 & K9x2a4);
	assign K9x2a4 = (~(Yjdw84 & X0v2a4));
	assign D9x2a4 = (R9x2a4 & Y9x2a4);
	assign Y9x2a4 = (~(Apyw84 & S1v2a4));
	assign R9x2a4 = (~(C80x84 & Z1v2a4));
	assign P8x2a4 = (Fax2a4 & Max2a4);
	assign Max2a4 = (~(Itgw84 & U2v2a4));
	assign Fax2a4 = (~(Q6fw84 & B3v2a4));
	assign B8x2a4 = (Tax2a4 & Abx2a4);
	assign Abx2a4 = (Hbx2a4 & Obx2a4);
	assign Obx2a4 = (~(S2kw84 & K4v2a4));
	assign Hbx2a4 = (~(Agiw84 & R4v2a4));
	assign Tax2a4 = (~(C8g2a4 | Vbx2a4));
	assign Vbx2a4 = (Gxbw84 & F5v2a4);
	assign G7x2a4 = (~(Oaaw84 & M5v2a4));
	assign E6x2a4 = (~(Qp63a4[27] & T5v2a4));
	assign HADDR[26] = (~(Ccx2a4 & Jcx2a4));
	assign Jcx2a4 = (~(Ao63a4[25] & F1hx84));
	assign Ccx2a4 = (Qcx2a4 & Xcx2a4);
	assign Xcx2a4 = (Kxu2a4 | Nxax84);
	assign Nxax84 = (!W2zx84);
	assign W2zx84 = (~(Edx2a4 & Ldx2a4));
	assign Ldx2a4 = (~(W6aw84 & M7ix84));
	assign Edx2a4 = (Sdx2a4 & Zdx2a4);
	assign Zdx2a4 = (~(Tyu2a4 & Gex2a4));
	assign Gex2a4 = (~(Nex2a4 & Uex2a4));
	assign Uex2a4 = (Bfx2a4 & Ifx2a4);
	assign Ifx2a4 = (Pfx2a4 & Wfx2a4);
	assign Wfx2a4 = (~(X0v2a4 & Cidw84));
	assign Pfx2a4 = (Dgx2a4 & Kgx2a4);
	assign Kgx2a4 = (~(S1v2a4 & Enyw84));
	assign Dgx2a4 = (~(Z1v2a4 & G60x84));
	assign Bfx2a4 = (Rgx2a4 & Ygx2a4);
	assign Ygx2a4 = (~(U2v2a4 & Mrgw84));
	assign Rgx2a4 = (~(B3v2a4 & U4fw84));
	assign Nex2a4 = (Fhx2a4 & Mhx2a4);
	assign Mhx2a4 = (Thx2a4 & Aix2a4);
	assign Aix2a4 = (~(K4v2a4 & W0kw84));
	assign Thx2a4 = (~(R4v2a4 & Eeiw84));
	assign Fhx2a4 = (~(H7g2a4 | Hix2a4));
	assign Hix2a4 = (F5v2a4 & Kvbw84);
	assign Sdx2a4 = (~(M5v2a4 & S8aw84));
	assign Qcx2a4 = (~(Qp63a4[26] & T5v2a4));
	assign HADDR[25] = (~(Oix2a4 & Vix2a4));
	assign Vix2a4 = (~(Ao63a4[24] & F1hx84));
	assign Oix2a4 = (Cjx2a4 & Jjx2a4);
	assign Jjx2a4 = (Kxu2a4 | Uxax84);
	assign Uxax84 = (!Dwyx84);
	assign Dwyx84 = (~(Qjx2a4 & Xjx2a4));
	assign Xjx2a4 = (~(A5aw84 & M7ix84));
	assign Qjx2a4 = (Ekx2a4 & Lkx2a4);
	assign Lkx2a4 = (~(Tyu2a4 & Skx2a4));
	assign Skx2a4 = (~(Zkx2a4 & Glx2a4));
	assign Glx2a4 = (Nlx2a4 & Ulx2a4);
	assign Ulx2a4 = (Bmx2a4 & Imx2a4);
	assign Imx2a4 = (~(Ggdw84 & X0v2a4));
	assign Bmx2a4 = (Pmx2a4 & Wmx2a4);
	assign Wmx2a4 = (~(Ilyw84 & S1v2a4));
	assign Pmx2a4 = (~(K40x84 & Z1v2a4));
	assign Nlx2a4 = (Dnx2a4 & Knx2a4);
	assign Knx2a4 = (~(Qpgw84 & U2v2a4));
	assign Dnx2a4 = (~(Y2fw84 & B3v2a4));
	assign Zkx2a4 = (Rnx2a4 & Ynx2a4);
	assign Ynx2a4 = (Fox2a4 & Mox2a4);
	assign Mox2a4 = (~(Azjw84 & K4v2a4));
	assign Fox2a4 = (~(Iciw84 & R4v2a4));
	assign Rnx2a4 = (~(J8g2a4 | Tox2a4));
	assign Tox2a4 = (Otbw84 & F5v2a4);
	assign Ekx2a4 = (~(W6aw84 & M5v2a4));
	assign Cjx2a4 = (~(Qp63a4[25] & T5v2a4));
	assign HADDR[24] = (~(Apx2a4 & Hpx2a4));
	assign Hpx2a4 = (~(Ao63a4[23] & F1hx84));
	assign Apx2a4 = (Opx2a4 & Vpx2a4);
	assign Vpx2a4 = (Kxu2a4 | Byax84);
	assign Byax84 = (!Tg1y84);
	assign Tg1y84 = (~(Cqx2a4 & Jqx2a4));
	assign Jqx2a4 = (~(E3aw84 & M7ix84));
	assign Cqx2a4 = (Qqx2a4 & Xqx2a4);
	assign Xqx2a4 = (~(Tyu2a4 & Erx2a4));
	assign Erx2a4 = (~(Lrx2a4 & Srx2a4));
	assign Srx2a4 = (Zrx2a4 & Gsx2a4);
	assign Gsx2a4 = (Nsx2a4 & Usx2a4);
	assign Usx2a4 = (~(Kedw84 & X0v2a4));
	assign Nsx2a4 = (Btx2a4 & Itx2a4);
	assign Itx2a4 = (~(Mjyw84 & S1v2a4));
	assign Btx2a4 = (~(O20x84 & Z1v2a4));
	assign Zrx2a4 = (Ptx2a4 & Wtx2a4);
	assign Wtx2a4 = (~(Ungw84 & U2v2a4));
	assign Ptx2a4 = (~(C1fw84 & B3v2a4));
	assign Lrx2a4 = (Dux2a4 & Kux2a4);
	assign Kux2a4 = (Rux2a4 & Yux2a4);
	assign Yux2a4 = (~(Exjw84 & K4v2a4));
	assign Rux2a4 = (~(Maiw84 & R4v2a4));
	assign Dux2a4 = (~(Lng2a4 | Fvx2a4));
	assign Fvx2a4 = (Srbw84 & F5v2a4);
	assign Qqx2a4 = (~(A5aw84 & M5v2a4));
	assign Opx2a4 = (~(T5v2a4 & Qp63a4[24]));
	assign HADDR[23] = (~(Mvx2a4 & Tvx2a4));
	assign Tvx2a4 = (~(Ao63a4[22] & F1hx84));
	assign Mvx2a4 = (Awx2a4 & Hwx2a4);
	assign Hwx2a4 = (Kxu2a4 | Iyax84);
	assign Iyax84 = (!L0zx84);
	assign L0zx84 = (~(Owx2a4 & Vwx2a4));
	assign Vwx2a4 = (~(I1aw84 & M7ix84));
	assign Owx2a4 = (Cxx2a4 & Jxx2a4);
	assign Jxx2a4 = (~(Tyu2a4 & Qxx2a4));
	assign Qxx2a4 = (~(Xxx2a4 & Eyx2a4));
	assign Eyx2a4 = (Lyx2a4 & Syx2a4);
	assign Syx2a4 = (Zyx2a4 & Gzx2a4);
	assign Gzx2a4 = (~(Ocdw84 & X0v2a4));
	assign Zyx2a4 = (Nzx2a4 & Uzx2a4);
	assign Uzx2a4 = (~(Qhyw84 & S1v2a4));
	assign Nzx2a4 = (~(S00x84 & Z1v2a4));
	assign Lyx2a4 = (B0y2a4 & I0y2a4);
	assign I0y2a4 = (~(Ylgw84 & U2v2a4));
	assign B0y2a4 = (~(Gzew84 & B3v2a4));
	assign Xxx2a4 = (P0y2a4 & W0y2a4);
	assign W0y2a4 = (D1y2a4 & K1y2a4);
	assign K1y2a4 = (~(Ivjw84 & K4v2a4));
	assign D1y2a4 = (~(Q8iw84 & R4v2a4));
	assign P0y2a4 = (~(Nog2a4 | R1y2a4));
	assign R1y2a4 = (Wpbw84 & F5v2a4);
	assign Cxx2a4 = (~(E3aw84 & M5v2a4));
	assign Awx2a4 = (~(Qp63a4[23] & T5v2a4));
	assign HADDR[22] = (~(Y1y2a4 & F2y2a4));
	assign F2y2a4 = (~(Ao63a4[21] & F1hx84));
	assign Y1y2a4 = (M2y2a4 & T2y2a4);
	assign T2y2a4 = (Kxu2a4 | Pyax84);
	assign Pyax84 = (!Xzyx84);
	assign Xzyx84 = (~(A3y2a4 & H3y2a4));
	assign H3y2a4 = (~(Mz9w84 & M7ix84));
	assign A3y2a4 = (O3y2a4 & V3y2a4);
	assign V3y2a4 = (~(Tyu2a4 & C4y2a4));
	assign C4y2a4 = (~(J4y2a4 & Q4y2a4));
	assign Q4y2a4 = (X4y2a4 & E5y2a4);
	assign E5y2a4 = (L5y2a4 & S5y2a4);
	assign S5y2a4 = (~(Sadw84 & X0v2a4));
	assign L5y2a4 = (Z5y2a4 & G6y2a4);
	assign G6y2a4 = (~(Ufyw84 & S1v2a4));
	assign Z5y2a4 = (~(Wyzw84 & Z1v2a4));
	assign X4y2a4 = (N6y2a4 & U6y2a4);
	assign U6y2a4 = (~(Ckgw84 & U2v2a4));
	assign N6y2a4 = (~(Kxew84 & B3v2a4));
	assign J4y2a4 = (B7y2a4 & I7y2a4);
	assign I7y2a4 = (P7y2a4 & W7y2a4);
	assign W7y2a4 = (~(Mtjw84 & K4v2a4));
	assign P7y2a4 = (~(U6iw84 & R4v2a4));
	assign B7y2a4 = (~(Sng2a4 | D8y2a4));
	assign D8y2a4 = (Aobw84 & F5v2a4);
	assign O3y2a4 = (~(I1aw84 & M5v2a4));
	assign M2y2a4 = (~(Qp63a4[22] & T5v2a4));
	assign HADDR[21] = (~(K8y2a4 & R8y2a4));
	assign R8y2a4 = (~(Ao63a4[20] & F1hx84));
	assign K8y2a4 = (Y8y2a4 & F9y2a4);
	assign F9y2a4 = (Kxu2a4 | Wyax84);
	assign Wyax84 = (!I2zx84);
	assign I2zx84 = (~(M9y2a4 & T9y2a4));
	assign T9y2a4 = (~(Qx9w84 & M7ix84));
	assign M9y2a4 = (Aay2a4 & Hay2a4);
	assign Hay2a4 = (~(Tyu2a4 & Oay2a4));
	assign Oay2a4 = (~(Vay2a4 & Cby2a4));
	assign Cby2a4 = (Jby2a4 & Qby2a4);
	assign Qby2a4 = (Xby2a4 & Ecy2a4);
	assign Ecy2a4 = (~(W8dw84 & X0v2a4));
	assign Xby2a4 = (Lcy2a4 & Scy2a4);
	assign Scy2a4 = (~(Ydyw84 & S1v2a4));
	assign Lcy2a4 = (~(Axzw84 & Z1v2a4));
	assign Jby2a4 = (Zcy2a4 & Gdy2a4);
	assign Gdy2a4 = (~(Gigw84 & U2v2a4));
	assign Zcy2a4 = (~(Ovew84 & B3v2a4));
	assign Vay2a4 = (Ndy2a4 & Udy2a4);
	assign Udy2a4 = (Bey2a4 & Iey2a4);
	assign Iey2a4 = (~(Qrjw84 & K4v2a4));
	assign Bey2a4 = (~(Y4iw84 & R4v2a4));
	assign Ndy2a4 = (~(Uog2a4 | Pey2a4));
	assign Pey2a4 = (Embw84 & F5v2a4);
	assign Aay2a4 = (~(Mz9w84 & M5v2a4));
	assign Y8y2a4 = (~(Qp63a4[21] & T5v2a4));
	assign HADDR[20] = (~(Wey2a4 & Dfy2a4));
	assign Dfy2a4 = (~(Ao63a4[19] & F1hx84));
	assign Wey2a4 = (Kfy2a4 & Rfy2a4);
	assign Rfy2a4 = (Kxu2a4 | Dzax84);
	assign Dzax84 = (!F4zx84);
	assign F4zx84 = (~(Yfy2a4 & Fgy2a4));
	assign Fgy2a4 = (~(Uv9w84 & M7ix84));
	assign Yfy2a4 = (Mgy2a4 & Tgy2a4);
	assign Tgy2a4 = (~(Tyu2a4 & Ahy2a4));
	assign Ahy2a4 = (~(Hhy2a4 & Ohy2a4));
	assign Ohy2a4 = (Vhy2a4 & Ciy2a4);
	assign Ciy2a4 = (Jiy2a4 & Qiy2a4);
	assign Qiy2a4 = (~(A7dw84 & X0v2a4));
	assign Jiy2a4 = (Xiy2a4 & Ejy2a4);
	assign Ejy2a4 = (~(Ccyw84 & S1v2a4));
	assign Xiy2a4 = (~(Evzw84 & Z1v2a4));
	assign Vhy2a4 = (Ljy2a4 & Sjy2a4);
	assign Sjy2a4 = (~(Kggw84 & U2v2a4));
	assign Ljy2a4 = (~(Stew84 & B3v2a4));
	assign Hhy2a4 = (Zjy2a4 & Gky2a4);
	assign Gky2a4 = (Nky2a4 & Uky2a4);
	assign Uky2a4 = (~(Upjw84 & K4v2a4));
	assign Nky2a4 = (~(C3iw84 & R4v2a4));
	assign Zjy2a4 = (~(Tkg2a4 | Bly2a4));
	assign Bly2a4 = (Ikbw84 & F5v2a4);
	assign Mgy2a4 = (~(Qx9w84 & M5v2a4));
	assign Kfy2a4 = (~(Qp63a4[20] & T5v2a4));
	assign HADDR[1] = (Xmu2a4 & Oya2a4);
	assign Oya2a4 = (~(Ily2a4 & Ply2a4));
	assign Ply2a4 = (~(T5v2a4 & Qp63a4[1]));
	assign Ily2a4 = (Wly2a4 & Dmy2a4);
	assign Dmy2a4 = (~(F1hx84 & Kmy2a4));
	assign Kmy2a4 = (~(Bzgx84 ^ Prax84));
	assign Wly2a4 = (Kxu2a4 | Kzax84);
	assign Kzax84 = (!Oi0y84);
	assign Oi0y84 = (~(Rmy2a4 & Ymy2a4));
	assign Ymy2a4 = (~(Cx8w84 & M7ix84));
	assign Rmy2a4 = (Fny2a4 & Mny2a4);
	assign Mny2a4 = (~(Tyu2a4 & Tny2a4));
	assign Tny2a4 = (~(Aoy2a4 & Hoy2a4));
	assign Hoy2a4 = (Ooy2a4 & Voy2a4);
	assign Voy2a4 = (Cpy2a4 & Jpy2a4);
	assign Jpy2a4 = (~(X0v2a4 & H8cw84));
	assign Cpy2a4 = (~(U2v2a4 & Rhfw84));
	assign Ooy2a4 = (Qpy2a4 & Xpy2a4);
	assign Xpy2a4 = (~(B3v2a4 & Zudw84));
	assign Qpy2a4 = (~(K4v2a4 & Briw84));
	assign Aoy2a4 = (~(Eqy2a4 | Evf2a4));
	assign Eqy2a4 = (~(Lqy2a4 & Sqy2a4));
	assign Sqy2a4 = (~(R4v2a4 & J4hw84));
	assign Lqy2a4 = (~(F5v2a4 & Plaw84));
	assign Fny2a4 = (~(M5v2a4 & Xy8w84));
	assign HADDR[19] = (~(Zqy2a4 & Gry2a4));
	assign Gry2a4 = (~(Ao63a4[18] & F1hx84));
	assign Zqy2a4 = (Nry2a4 & Ury2a4);
	assign Ury2a4 = (Kxu2a4 | Rzax84);
	assign Rzax84 = (!Yu0y84);
	assign Yu0y84 = (~(Bsy2a4 & Isy2a4));
	assign Isy2a4 = (~(Yt9w84 & M7ix84));
	assign Bsy2a4 = (Psy2a4 & Wsy2a4);
	assign Wsy2a4 = (~(Tyu2a4 & Dty2a4));
	assign Dty2a4 = (~(Kty2a4 & Rty2a4));
	assign Rty2a4 = (Yty2a4 & Fuy2a4);
	assign Fuy2a4 = (Muy2a4 & Tuy2a4);
	assign Tuy2a4 = (~(E5dw84 & X0v2a4));
	assign Muy2a4 = (Avy2a4 & Hvy2a4);
	assign Hvy2a4 = (~(Gayw84 & S1v2a4));
	assign Avy2a4 = (~(Itzw84 & Z1v2a4));
	assign Yty2a4 = (Ovy2a4 & Vvy2a4);
	assign Vvy2a4 = (~(Oegw84 & U2v2a4));
	assign Ovy2a4 = (~(Wrew84 & B3v2a4));
	assign Kty2a4 = (Cwy2a4 & Jwy2a4);
	assign Jwy2a4 = (Qwy2a4 & Xwy2a4);
	assign Xwy2a4 = (~(Ynjw84 & K4v2a4));
	assign Qwy2a4 = (~(G1iw84 & R4v2a4));
	assign Cwy2a4 = (~(Vlg2a4 | Exy2a4));
	assign Exy2a4 = (Mibw84 & F5v2a4);
	assign Psy2a4 = (~(Uv9w84 & M5v2a4));
	assign Nry2a4 = (~(T5v2a4 & Qp63a4[19]));
	assign HADDR[18] = (~(Lxy2a4 & Sxy2a4));
	assign Sxy2a4 = (~(Ao63a4[17] & F1hx84));
	assign Lxy2a4 = (Zxy2a4 & Gyy2a4);
	assign Gyy2a4 = (Kxu2a4 | Yzax84);
	assign Yzax84 = (!Ns0y84);
	assign Ns0y84 = (~(Nyy2a4 & Uyy2a4));
	assign Uyy2a4 = (~(Cs9w84 & M7ix84));
	assign Nyy2a4 = (Bzy2a4 & Izy2a4);
	assign Izy2a4 = (~(Tyu2a4 & Pzy2a4));
	assign Pzy2a4 = (~(Wzy2a4 & D0z2a4));
	assign D0z2a4 = (K0z2a4 & R0z2a4);
	assign R0z2a4 = (Y0z2a4 & F1z2a4);
	assign F1z2a4 = (~(I3dw84 & X0v2a4));
	assign Y0z2a4 = (M1z2a4 & T1z2a4);
	assign T1z2a4 = (~(K8yw84 & S1v2a4));
	assign M1z2a4 = (~(Mrzw84 & Z1v2a4));
	assign K0z2a4 = (A2z2a4 & H2z2a4);
	assign H2z2a4 = (~(Scgw84 & U2v2a4));
	assign A2z2a4 = (~(Aqew84 & B3v2a4));
	assign Wzy2a4 = (O2z2a4 & V2z2a4);
	assign V2z2a4 = (C3z2a4 & J3z2a4);
	assign J3z2a4 = (~(Cmjw84 & K4v2a4));
	assign C3z2a4 = (~(Kzhw84 & R4v2a4));
	assign O2z2a4 = (~(Alg2a4 | Q3z2a4));
	assign Q3z2a4 = (Qgbw84 & F5v2a4);
	assign Bzy2a4 = (~(Yt9w84 & M5v2a4));
	assign Zxy2a4 = (~(T5v2a4 & Qp63a4[18]));
	assign HADDR[17] = (~(X3z2a4 & E4z2a4));
	assign E4z2a4 = (~(Ao63a4[16] & F1hx84));
	assign X3z2a4 = (L4z2a4 & S4z2a4);
	assign S4z2a4 = (Kxu2a4 | F0bx84);
	assign F0bx84 = (!Ie1y84);
	assign Ie1y84 = (~(Z4z2a4 & G5z2a4));
	assign G5z2a4 = (~(Gq9w84 & M7ix84));
	assign Z4z2a4 = (N5z2a4 & U5z2a4);
	assign U5z2a4 = (~(Tyu2a4 & B6z2a4));
	assign B6z2a4 = (~(I6z2a4 & P6z2a4));
	assign P6z2a4 = (W6z2a4 & D7z2a4);
	assign D7z2a4 = (K7z2a4 & R7z2a4);
	assign R7z2a4 = (~(M1dw84 & X0v2a4));
	assign K7z2a4 = (Y7z2a4 & F8z2a4);
	assign F8z2a4 = (~(O6yw84 & S1v2a4));
	assign Y7z2a4 = (~(Qpzw84 & Z1v2a4));
	assign W6z2a4 = (M8z2a4 & T8z2a4);
	assign T8z2a4 = (~(Wagw84 & U2v2a4));
	assign M8z2a4 = (~(Eoew84 & B3v2a4));
	assign I6z2a4 = (A9z2a4 & H9z2a4);
	assign H9z2a4 = (O9z2a4 & V9z2a4);
	assign V9z2a4 = (~(Gkjw84 & K4v2a4));
	assign O9z2a4 = (~(Oxhw84 & R4v2a4));
	assign A9z2a4 = (~(Cmg2a4 | Caz2a4));
	assign Caz2a4 = (Uebw84 & F5v2a4);
	assign N5z2a4 = (~(Cs9w84 & M5v2a4));
	assign L4z2a4 = (~(T5v2a4 & Qp63a4[17]));
	assign HADDR[16] = (~(Jaz2a4 & Qaz2a4));
	assign Qaz2a4 = (~(Ao63a4[15] & F1hx84));
	assign Jaz2a4 = (Xaz2a4 & Ebz2a4);
	assign Ebz2a4 = (Kxu2a4 | M0bx84);
	assign M0bx84 = (!K3zx84);
	assign K3zx84 = (~(Lbz2a4 & Sbz2a4));
	assign Sbz2a4 = (~(Ko9w84 & M7ix84));
	assign Lbz2a4 = (Zbz2a4 & Gcz2a4);
	assign Gcz2a4 = (~(Tyu2a4 & Ncz2a4));
	assign Ncz2a4 = (~(Ucz2a4 & Bdz2a4));
	assign Bdz2a4 = (Idz2a4 & Pdz2a4);
	assign Pdz2a4 = (Wdz2a4 & Dez2a4);
	assign Dez2a4 = (~(Qzcw84 & X0v2a4));
	assign Wdz2a4 = (Kez2a4 & Rez2a4);
	assign Rez2a4 = (~(S4yw84 & S1v2a4));
	assign Kez2a4 = (~(Unzw84 & Z1v2a4));
	assign Idz2a4 = (Yez2a4 & Ffz2a4);
	assign Ffz2a4 = (~(A9gw84 & U2v2a4));
	assign Yez2a4 = (~(Imew84 & B3v2a4));
	assign Ucz2a4 = (Mfz2a4 & Tfz2a4);
	assign Tfz2a4 = (Agz2a4 & Hgz2a4);
	assign Hgz2a4 = (~(Kijw84 & K4v2a4));
	assign Agz2a4 = (~(Svhw84 & R4v2a4));
	assign Mfz2a4 = (~(Oeg2a4 | Ogz2a4));
	assign Ogz2a4 = (Ycbw84 & F5v2a4);
	assign Zbz2a4 = (~(Gq9w84 & M5v2a4));
	assign Xaz2a4 = (~(Qp63a4[16] & T5v2a4));
	assign HADDR[15] = (~(Vgz2a4 & Chz2a4));
	assign Chz2a4 = (~(Ao63a4[14] & F1hx84));
	assign Vgz2a4 = (Jhz2a4 & Qhz2a4);
	assign Qhz2a4 = (Kxu2a4 | T0bx84);
	assign T0bx84 = (!Bvyx84);
	assign Bvyx84 = (~(Xhz2a4 & Eiz2a4));
	assign Eiz2a4 = (~(Om9w84 & M7ix84));
	assign Xhz2a4 = (Liz2a4 & Siz2a4);
	assign Siz2a4 = (~(Tyu2a4 & Ziz2a4));
	assign Ziz2a4 = (~(Gjz2a4 & Njz2a4));
	assign Njz2a4 = (Ujz2a4 & Bkz2a4);
	assign Bkz2a4 = (Ikz2a4 & Pkz2a4);
	assign Pkz2a4 = (~(X0v2a4 & Uxcw84));
	assign Ikz2a4 = (Wkz2a4 & Dlz2a4);
	assign Dlz2a4 = (~(S1v2a4 & W2yw84));
	assign Wkz2a4 = (~(Z1v2a4 & Ylzw84));
	assign Ujz2a4 = (Klz2a4 & Rlz2a4);
	assign Rlz2a4 = (~(U2v2a4 & E7gw84));
	assign Klz2a4 = (~(B3v2a4 & Mkew84));
	assign Gjz2a4 = (Ylz2a4 & Fmz2a4);
	assign Fmz2a4 = (Mmz2a4 & Tmz2a4);
	assign Tmz2a4 = (~(K4v2a4 & Ogjw84));
	assign Mmz2a4 = (~(R4v2a4 & Wthw84));
	assign Ylz2a4 = (~(Qfg2a4 | Anz2a4));
	assign Anz2a4 = (F5v2a4 & Cbbw84);
	assign Liz2a4 = (~(M5v2a4 & Ko9w84));
	assign Jhz2a4 = (~(Qp63a4[15] & T5v2a4));
	assign HADDR[14] = (~(Hnz2a4 & Onz2a4));
	assign Onz2a4 = (~(Ao63a4[13] & F1hx84));
	assign Hnz2a4 = (Vnz2a4 & Coz2a4);
	assign Coz2a4 = (Kxu2a4 | A1bx84);
	assign A1bx84 = (!Vyyx84);
	assign Vyyx84 = (~(Joz2a4 & Qoz2a4));
	assign Qoz2a4 = (~(Sk9w84 & M7ix84));
	assign Joz2a4 = (Xoz2a4 & Epz2a4);
	assign Epz2a4 = (~(Tyu2a4 & Lpz2a4));
	assign Lpz2a4 = (~(Spz2a4 & Zpz2a4));
	assign Zpz2a4 = (Gqz2a4 & Nqz2a4);
	assign Nqz2a4 = (Uqz2a4 & Brz2a4);
	assign Brz2a4 = (~(Yvcw84 & X0v2a4));
	assign Uqz2a4 = (Irz2a4 & Prz2a4);
	assign Prz2a4 = (~(A1yw84 & S1v2a4));
	assign Irz2a4 = (~(Ckzw84 & Z1v2a4));
	assign Gqz2a4 = (Wrz2a4 & Dsz2a4);
	assign Dsz2a4 = (~(I5gw84 & U2v2a4));
	assign Wrz2a4 = (~(Qiew84 & B3v2a4));
	assign Spz2a4 = (Ksz2a4 & Rsz2a4);
	assign Rsz2a4 = (Ysz2a4 & Ftz2a4);
	assign Ftz2a4 = (~(Sejw84 & K4v2a4));
	assign Ysz2a4 = (~(Ashw84 & R4v2a4));
	assign Ksz2a4 = (~(Veg2a4 | Mtz2a4));
	assign Mtz2a4 = (G9bw84 & F5v2a4);
	assign Xoz2a4 = (~(Om9w84 & M5v2a4));
	assign Vnz2a4 = (~(Qp63a4[14] & T5v2a4));
	assign HADDR[13] = (~(Ttz2a4 & Auz2a4));
	assign Auz2a4 = (~(Ao63a4[12] & F1hx84));
	assign Ttz2a4 = (Huz2a4 & Ouz2a4);
	assign Ouz2a4 = (Kxu2a4 | H1bx84);
	assign H1bx84 = (!Rwyx84);
	assign Rwyx84 = (~(Vuz2a4 & Cvz2a4));
	assign Cvz2a4 = (~(Wi9w84 & M7ix84));
	assign Vuz2a4 = (Jvz2a4 & Qvz2a4);
	assign Qvz2a4 = (~(Tyu2a4 & Xvz2a4));
	assign Xvz2a4 = (~(Ewz2a4 & Lwz2a4));
	assign Lwz2a4 = (Swz2a4 & Zwz2a4);
	assign Zwz2a4 = (Gxz2a4 & Nxz2a4);
	assign Nxz2a4 = (~(Cucw84 & X0v2a4));
	assign Gxz2a4 = (Uxz2a4 & Byz2a4);
	assign Byz2a4 = (~(Ezxw84 & S1v2a4));
	assign Uxz2a4 = (~(Gizw84 & Z1v2a4));
	assign Swz2a4 = (Iyz2a4 & Pyz2a4);
	assign Pyz2a4 = (~(M3gw84 & U2v2a4));
	assign Iyz2a4 = (~(Ugew84 & B3v2a4));
	assign Ewz2a4 = (Wyz2a4 & Dzz2a4);
	assign Dzz2a4 = (Kzz2a4 & Rzz2a4);
	assign Rzz2a4 = (~(Wcjw84 & K4v2a4));
	assign Kzz2a4 = (~(Eqhw84 & R4v2a4));
	assign Wyz2a4 = (~(Xfg2a4 | Yzz2a4));
	assign Yzz2a4 = (K7bw84 & F5v2a4);
	assign Jvz2a4 = (~(Sk9w84 & M5v2a4));
	assign Huz2a4 = (~(Qp63a4[13] & T5v2a4));
	assign HADDR[12] = (~(F003a4 & M003a4));
	assign M003a4 = (~(Ao63a4[11] & F1hx84));
	assign F003a4 = (T003a4 & A103a4);
	assign A103a4 = (Kxu2a4 | O1bx84);
	assign O1bx84 = (!W01y84);
	assign W01y84 = (~(H103a4 & O103a4));
	assign O103a4 = (~(Ah9w84 & M7ix84));
	assign H103a4 = (V103a4 & C203a4);
	assign C203a4 = (~(Tyu2a4 & J203a4));
	assign J203a4 = (~(Q203a4 & X203a4));
	assign X203a4 = (E303a4 & L303a4);
	assign L303a4 = (S303a4 & Z303a4);
	assign Z303a4 = (~(Gscw84 & X0v2a4));
	assign S303a4 = (G403a4 & N403a4);
	assign N403a4 = (~(Ixxw84 & S1v2a4));
	assign G403a4 = (~(Kgzw84 & Z1v2a4));
	assign E303a4 = (U403a4 & B503a4);
	assign B503a4 = (~(Q1gw84 & U2v2a4));
	assign U403a4 = (~(Yeew84 & B3v2a4));
	assign Q203a4 = (I503a4 & P503a4);
	assign P503a4 = (W503a4 & D603a4);
	assign D603a4 = (~(Abjw84 & K4v2a4));
	assign W503a4 = (~(Iohw84 & R4v2a4));
	assign I503a4 = (~(Wbg2a4 | K603a4));
	assign K603a4 = (O5bw84 & F5v2a4);
	assign V103a4 = (~(Wi9w84 & M5v2a4));
	assign T003a4 = (~(T5v2a4 & Qp63a4[12]));
	assign HADDR[11] = (~(R603a4 & Y603a4));
	assign Y603a4 = (~(Ao63a4[10] & F1hx84));
	assign R603a4 = (F703a4 & M703a4);
	assign M703a4 = (Kxu2a4 | V1bx84);
	assign V1bx84 = (!Txyx84);
	assign Txyx84 = (~(T703a4 & A803a4));
	assign A803a4 = (~(Ef9w84 & M7ix84));
	assign T703a4 = (H803a4 & O803a4);
	assign O803a4 = (~(Tyu2a4 & V803a4));
	assign V803a4 = (~(C903a4 & J903a4));
	assign J903a4 = (Q903a4 & X903a4);
	assign X903a4 = (Ea03a4 & La03a4);
	assign La03a4 = (~(Kqcw84 & X0v2a4));
	assign Ea03a4 = (Sa03a4 & Za03a4);
	assign Za03a4 = (~(Mvxw84 & S1v2a4));
	assign Sa03a4 = (~(Oezw84 & Z1v2a4));
	assign Q903a4 = (Gb03a4 & Nb03a4);
	assign Nb03a4 = (~(Uzfw84 & U2v2a4));
	assign Gb03a4 = (~(Cdew84 & B3v2a4));
	assign C903a4 = (Ub03a4 & Bc03a4);
	assign Bc03a4 = (Ic03a4 & Pc03a4);
	assign Pc03a4 = (~(E9jw84 & K4v2a4));
	assign Ic03a4 = (~(Mmhw84 & R4v2a4));
	assign Ub03a4 = (~(Ycg2a4 | Wc03a4));
	assign Wc03a4 = (S3bw84 & F5v2a4);
	assign H803a4 = (~(Ah9w84 & M5v2a4));
	assign F703a4 = (~(Qp63a4[11] & T5v2a4));
	assign HADDR[10] = (~(Dd03a4 & Kd03a4));
	assign Kd03a4 = (~(Ao63a4[9] & F1hx84));
	assign F1hx84 = (!Dkix84);
	assign Dd03a4 = (Rd03a4 & Yd03a4);
	assign Yd03a4 = (Kxu2a4 | C2bx84);
	assign C2bx84 = (!Fxyx84);
	assign Fxyx84 = (~(Fe03a4 & Me03a4));
	assign Me03a4 = (~(Jd9w84 & M7ix84));
	assign Fe03a4 = (Te03a4 & Af03a4);
	assign Af03a4 = (~(Tyu2a4 & Hf03a4));
	assign Hf03a4 = (~(Of03a4 & Vf03a4));
	assign Vf03a4 = (Cg03a4 & Jg03a4);
	assign Jg03a4 = (Qg03a4 & Xg03a4);
	assign Xg03a4 = (~(Oocw84 & X0v2a4));
	assign Qg03a4 = (Eh03a4 & Lh03a4);
	assign Lh03a4 = (~(Qtxw84 & S1v2a4));
	assign S1v2a4 = (Sh03a4 & Zh03a4);
	assign Sh03a4 = (Gi03a4 & Mdxw84);
	assign Eh03a4 = (~(Sczw84 & Z1v2a4));
	assign Z1v2a4 = (Ni03a4 & Zh03a4);
	assign Ni03a4 = (Gi03a4 & Fvfx84);
	assign Fvfx84 = (!Mdxw84);
	assign Cg03a4 = (Ui03a4 & Bj03a4);
	assign Bj03a4 = (~(Yxfw84 & U2v2a4));
	assign Ui03a4 = (~(Gbew84 & B3v2a4));
	assign Of03a4 = (Ij03a4 & Pj03a4);
	assign Pj03a4 = (Wj03a4 & Dk03a4);
	assign Dk03a4 = (~(I7jw84 & K4v2a4));
	assign Wj03a4 = (~(Qkhw84 & R4v2a4));
	assign Ij03a4 = (~(Dcg2a4 | Kk03a4));
	assign Kk03a4 = (W1bw84 & F5v2a4);
	assign Te03a4 = (~(Ef9w84 & M5v2a4));
	assign Rd03a4 = (~(Qp63a4[10] & T5v2a4));
	assign HADDR[0] = (Rk03a4 & Xmu2a4);
	assign Xmu2a4 = (N6r2a4 & Alu2a4);
	assign Alu2a4 = (~(Yk03a4 & O2hx84));
	assign O2hx84 = (Fl03a4 & Ml03a4);
	assign Ml03a4 = (Tl03a4 & Am03a4);
	assign Am03a4 = (Hm03a4 & Om03a4);
	assign Om03a4 = (Vm03a4 & Rsl2a4);
	assign Rsl2a4 = (~(Cn03a4 & Zvix84));
	assign Zvix84 = (Zo2x84 & Bw2x84);
	assign Cn03a4 = (~(H6dx84 | Jnix84));
	assign Vm03a4 = (~(Jn03a4 & Gwix84));
	assign Jn03a4 = (~(Wbcx84 | Ewax84));
	assign Wbcx84 = (!Wlnx84);
	assign Hm03a4 = (Qn03a4 & Xn03a4);
	assign Xn03a4 = (~(N4ix84 & Eo03a4));
	assign Eo03a4 = (~(Lo03a4 & So03a4));
	assign So03a4 = (Zo03a4 & Gp03a4);
	assign Gp03a4 = (~(Np03a4 & Aq42a4));
	assign Np03a4 = (~(Ewax84 | D4dx84));
	assign Zo03a4 = (~(Up03a4 | Bf52a4));
	assign Bf52a4 = (Soix84 & Ambx84);
	assign Up03a4 = (Bq03a4 & E3ix84);
	assign Bq03a4 = (~(Ambx84 | Yrbx84));
	assign Yrbx84 = (!Vzcx84);
	assign Lo03a4 = (Iq03a4 & Pq03a4);
	assign Pq03a4 = (~(Y1gx84 & F2gx84));
	assign Iq03a4 = (Qhl2a4 & Wq03a4);
	assign Wq03a4 = (~(Pxbx84 & Dr03a4));
	assign Dr03a4 = (~(Hkdx84 & Kr03a4));
	assign Kr03a4 = (~(Laix84 & Drbx84));
	assign Laix84 = (Tsix84 & Ewax84);
	assign Hkdx84 = (!Ozcx84);
	assign Qhl2a4 = (V2ox84 | Hu2x84);
	assign V2ox84 = (!Afix84);
	assign Afix84 = (Fn2x84 & Rvlx84);
	assign Qn03a4 = (~(Rr03a4 & Nacx84));
	assign Rr03a4 = (~(Mg62a4 | Hu2x84));
	assign Mg62a4 = (!Zymx84);
	assign Tl03a4 = (Yr03a4 & Fs03a4);
	assign Fs03a4 = (~(Ms03a4 & F2gx84));
	assign Ms03a4 = (Ts03a4 & Gpbx84);
	assign Ts03a4 = (~(At03a4 & Ht03a4));
	assign Ht03a4 = (B5bx84 | Ns2x84);
	assign At03a4 = (Fycx84 | D4dx84);
	assign Yr03a4 = (Ot03a4 & Vt03a4);
	assign Vt03a4 = (~(Ffox84 & Mmvx84));
	assign Ot03a4 = (~(Cu03a4 & Uwix84));
	assign Cu03a4 = (~(Ambx84 | Ns2x84));
	assign Fl03a4 = (Ju03a4 & Qu03a4);
	assign Qu03a4 = (Xu03a4 & Ev03a4);
	assign Ev03a4 = (Lv03a4 & Jxfx84);
	assign Jxfx84 = (~(Yzhx84 & A7cx84));
	assign Lv03a4 = (~(Sv03a4 & Cavx84));
	assign Cavx84 = (Tq2x84 & Qxmx84);
	assign Sv03a4 = (~(Lrfx84 | Zo2x84));
	assign Lrfx84 = (!Rvlx84);
	assign Xu03a4 = (Zv03a4 & Gw03a4);
	assign Gw03a4 = (~(Nw03a4 & Uw03a4));
	assign Uw03a4 = (~(Kd82a4 | Klvx84));
	assign Klvx84 = (Gz4w84 & Ns2x84);
	assign Kd82a4 = (Hu2x84 & Ns2x84);
	assign Nw03a4 = (Bx03a4 & Pz2x84);
	assign Bx03a4 = (Wqbx84 ? Ix03a4 : Vnl2a4);
	assign Zv03a4 = (~(Px03a4 & Ix03a4));
	assign Ix03a4 = (Wx03a4 & Pxbx84);
	assign Wx03a4 = (~(Hgvx84 | Mmvx84));
	assign Px03a4 = (~(Tsix84 | Yybx84));
	assign Yybx84 = (!Fg62a4);
	assign Fg62a4 = (~(Dy03a4 & Ky03a4));
	assign Ky03a4 = (Ry03a4 & Tk63a4[27]);
	assign Ry03a4 = (Bg5w84 & W7gx84);
	assign W7gx84 = (~(Yy03a4 & Wcm2a4));
	assign Wcm2a4 = (Icm2a4 & K7e2a4);
	assign K7e2a4 = (!Nj63a4[3]);
	assign Icm2a4 = (~(Nj63a4[4] | Nj63a4[5]));
	assign Yy03a4 = (Fz03a4 & Tbb2a4);
	assign Tbb2a4 = (!Nj63a4[0]);
	assign Fz03a4 = (~(Nj63a4[1] | Nj63a4[2]));
	assign Dy03a4 = (Mz03a4 & Tk63a4[30]);
	assign Mz03a4 = (Tk63a4[29] & Tk63a4[28]);
	assign Ju03a4 = (Tz03a4 & Dccx84);
	assign Tz03a4 = (A013a4 & H013a4);
	assign H013a4 = (~(O013a4 & G4wx84));
	assign G4wx84 = (N052a4 & Vzcx84);
	assign N052a4 = (V013a4 & Tk63a4[2]);
	assign V013a4 = (Lo4w84 & We62a4);
	assign We62a4 = (!Ws4w84);
	assign O013a4 = (~(Yrix84 | Ambx84));
	assign A013a4 = (O2ox84 | Rmnx84);
	assign Rmnx84 = (!Uj2x84);
	assign Yk03a4 = (C113a4 & J113a4);
	assign J113a4 = (~(Q113a4 & X113a4));
	assign X113a4 = (~(E213a4 & Gz4w84));
	assign E213a4 = (~(Ya2x84 | Ih0x84));
	assign Q113a4 = (~(L213a4 & S213a4));
	assign S213a4 = (Bzgx84 | Jrlx84);
	assign Jrlx84 = (!Dsax84);
	assign Dsax84 = (Bi2x84 & Z213a4);
	assign L213a4 = (Tplx84 | Aqlx84);
	assign Tplx84 = (~(Soix84 & Mnux84));
	assign Soix84 = (Jm92a4 & Zgxx84);
	assign Jm92a4 = (Gpbx84 & G4bx84);
	assign C113a4 = (~(Prax84 & Bzgx84));
	assign Bzgx84 = (!Tk63a4[0]);
	assign Prax84 = (Ig2x84 & Z213a4);
	assign Z213a4 = (!Aqlx84);
	assign Aqlx84 = (~(Fnux84 | G313a4));
	assign G313a4 = (!Mnux84);
	assign Mnux84 = (~(N313a4 & U313a4));
	assign U313a4 = (B413a4 & I413a4);
	assign I413a4 = (P413a4 & W413a4);
	assign W413a4 = (~(D513a4 & J982a4));
	assign D513a4 = (Y3i2a4 & Vx2x84);
	assign P413a4 = (~(V4c2a4 | Qn82a4));
	assign Qn82a4 = (Rvlx84 & Vx2x84);
	assign Rvlx84 = (J13x84 & Bw2x84);
	assign V4c2a4 = (Zoix84 & Wlnx84);
	assign Zoix84 = (~(Xcmx84 | Tswx84));
	assign Xcmx84 = (!D9mx84);
	assign B413a4 = (K513a4 & R513a4);
	assign R513a4 = (~(Y513a4 & H6dx84));
	assign Y513a4 = (~(F613a4 & M613a4));
	assign M613a4 = (~(T613a4 & On72a4));
	assign F613a4 = (A713a4 & H713a4);
	assign H713a4 = (~(O713a4 & Zymx84));
	assign Zymx84 = (N4ix84 & Ambx84);
	assign O713a4 = (~(Kzvx84 | Tq2x84));
	assign Kzvx84 = (B5bx84 | Yqcx84);
	assign A713a4 = (~(V713a4 & Sbvx84));
	assign V713a4 = (~(N4ix84 | Fn2x84));
	assign K513a4 = (C813a4 & J813a4);
	assign J813a4 = (~(Q0yx84 & J0dx84));
	assign J0dx84 = (~(Fthx84 | G4bx84));
	assign C813a4 = (Q813a4 | J13x84);
	assign N313a4 = (X813a4 & E913a4);
	assign E913a4 = (L913a4 & S913a4);
	assign S913a4 = (~(G33x84 & Z913a4));
	assign Z913a4 = (~(Ga13a4 & Na13a4));
	assign Na13a4 = (Ua13a4 & Bb13a4);
	assign Bb13a4 = (~(Ib13a4 & F7bx84));
	assign Ib13a4 = (Tamx84 & Pb13a4);
	assign Pb13a4 = (~(N4bx84 & Wb13a4));
	assign Wb13a4 = (B3dx84 | El42a4);
	assign El42a4 = (!Rv42a4);
	assign Rv42a4 = (~(Nrnx84 & Dc13a4));
	assign Dc13a4 = (Iicx84 | Jmcx84);
	assign Jmcx84 = (!Ey5w84);
	assign Iicx84 = (!Wz5w84);
	assign Nrnx84 = (O16w84 & Qzkx84);
	assign Qzkx84 = (!G36w84);
	assign B3dx84 = (!Deox84);
	assign N4bx84 = (!Yzhx84);
	assign Tamx84 = (~(Qtcx84 | Ub6w84));
	assign Qtcx84 = (!E8dx84);
	assign Ua13a4 = (~(Kc13a4 & Hwmx84));
	assign Hwmx84 = (~(P1mx84 | Fn2x84));
	assign P1mx84 = (!Nr62a4);
	assign Kc13a4 = (D9mx84 & Rc13a4);
	assign Rc13a4 = (~(Qcmx84 & Yc13a4));
	assign Yc13a4 = (T692a4 | W05w84);
	assign T692a4 = (Plnx84 | Tp42a4);
	assign Tp42a4 = (Gf6w84 & Oxlx84);
	assign Oxlx84 = (~(J8cx84 | Iokx84));
	assign Plnx84 = (C2ix84 & Iokx84);
	assign C2ix84 = (Zg6w84 & Xlkx84);
	assign Qcmx84 = (!Jtcx84);
	assign Ga13a4 = (Dccx84 & Fd13a4);
	assign Fd13a4 = (~(Md13a4 & Yqcx84));
	assign Md13a4 = (~(Td13a4 & Ae13a4));
	assign Ae13a4 = (~(F7bx84 & He13a4));
	assign He13a4 = (~(Oe13a4 & Ve13a4));
	assign Ve13a4 = (~(Edmx84 & Iokx84));
	assign Edmx84 = (~(Ouhx84 | J8cx84));
	assign Ouhx84 = (!Fhmx84);
	assign Fhmx84 = (Gf6w84 & Hgvx84);
	assign Oe13a4 = (~(Cf13a4 | Pcix84));
	assign Pcix84 = (Jtcx84 & Hgvx84);
	assign Jtcx84 = (Xlkx84 & J8cx84);
	assign J8cx84 = (!Zg6w84);
	assign Xlkx84 = (!Gf6w84);
	assign Cf13a4 = (E8dx84 & Jf13a4);
	assign Jf13a4 = (~(Zg6w84 & Qf13a4));
	assign Qf13a4 = (Iokx84 | Gf6w84);
	assign Iokx84 = (!Ub6w84);
	assign E8dx84 = (Hgvx84 & F3mx84);
	assign F3mx84 = (!W05w84);
	assign F7bx84 = (Vx2x84 & G4bx84);
	assign Td13a4 = (~(Y3i2a4 & F352a4));
	assign Dccx84 = (Xf13a4 & Ewl2a4);
	assign Ewl2a4 = (Axb2a4 | Tq2x84);
	assign Axb2a4 = (!Y0hx84);
	assign Y0hx84 = (D53x84 & Ambx84);
	assign Xf13a4 = (H6dx84 | Kxcx84);
	assign Kxcx84 = (!On72a4);
	assign L913a4 = (Eg13a4 & Lg13a4);
	assign Lg13a4 = (~(T0px84 & Sbvx84));
	assign T0px84 = (Livx84 & Mmvx84);
	assign Eg13a4 = (~(Atix84 & Sg13a4));
	assign Sg13a4 = (~(I2b2a4 & Zg13a4));
	assign Zg13a4 = (Gh13a4 & Nh13a4);
	assign Nh13a4 = (Yqcx84 | Tq2x84);
	assign Gh13a4 = (~(Uh13a4 | Vnl2a4));
	assign Vnl2a4 = (F2gx84 & Vx2x84);
	assign Uh13a4 = (~(Wqbx84 | Fn2x84));
	assign I2b2a4 = (~(Qxmx84 | Pqbx84));
	assign Atix84 = (Gz4w84 & H6dx84);
	assign X813a4 = (Bi13a4 & Ii13a4);
	assign Ii13a4 = (Undx84 ? Wi13a4 : Pi13a4);
	assign Wi13a4 = (~(Gwix84 & Dj13a4));
	assign Dj13a4 = (~(Evix84 & Kj13a4));
	assign Kj13a4 = (H6dx84 | Tsix84);
	assign Pi13a4 = (~(Nndx84 & Hgvx84));
	assign Nndx84 = (Wqbx84 & Pqbx84);
	assign Bi13a4 = (Rj13a4 & Yj13a4);
	assign Yj13a4 = (~(Y6bx84 & A7cx84));
	assign A7cx84 = (~(Ambx84 | Qxmx84));
	assign Rj13a4 = (~(P0gx84 & Hu2x84));
	assign P0gx84 = (Nr62a4 & Ambx84);
	assign Nr62a4 = (Bw2x84 & Wqbx84);
	assign Fnux84 = (!R3ex84);
	assign R3ex84 = (~(Fk13a4 & Mk13a4));
	assign Mk13a4 = (~(Y1gx84 & Pz2x84));
	assign Fk13a4 = (Tk13a4 & Iyl2a4);
	assign Iyl2a4 = (~(G52y84 & Y3i2a4));
	assign G52y84 = (~(Gz4w84 | Zo2x84));
	assign Tk13a4 = (~(Al13a4 & Mmvx84));
	assign Al13a4 = (~(Fthx84 & Hl13a4));
	assign Hl13a4 = (Rybx84 | D4dx84);
	assign Rybx84 = (!S3ix84);
	assign Rk03a4 = (~(Cza2a4 | Htt2a4));
	assign Htt2a4 = (!N1p2a4);
	assign N1p2a4 = (~(N6r2a4 & Ol13a4));
	assign Ol13a4 = (~(Vl13a4 & Cm13a4));
	assign Cm13a4 = (Ewax84 ? Dybx84 : S1dx84);
	assign Dybx84 = (!Lw72a4);
	assign Vl13a4 = (Jm13a4 & F5dx84);
	assign F5dx84 = (!J982a4);
	assign J982a4 = (Hu2x84 & Tq2x84);
	assign Jm13a4 = (Fycx84 | Ns2x84);
	assign N6r2a4 = (Qm13a4 & Xm13a4);
	assign Xm13a4 = (En13a4 & Ambx84);
	assign En13a4 = (Pqbx84 | Evix84);
	assign Qm13a4 = (~(Ln13a4 | Sq62a4));
	assign Sq62a4 = (Xm92a4 & Undx84);
	assign Ln13a4 = (~(H8px84 | On72a4));
	assign Cza2a4 = (Sn13a4 & Zn13a4);
	assign Zn13a4 = (Kxu2a4 | J2bx84);
	assign J2bx84 = (!Cq0y84);
	assign Cq0y84 = (~(Go13a4 & No13a4));
	assign No13a4 = (~(Tyu2a4 & Uo13a4));
	assign Uo13a4 = (~(Bp13a4 & Ip13a4));
	assign Ip13a4 = (Pp13a4 & Wp13a4);
	assign Wp13a4 = (Dq13a4 & Kq13a4);
	assign Kq13a4 = (~(X0v2a4 & M6cw84));
	assign X0v2a4 = (Rq13a4 & Gi03a4);
	assign Dq13a4 = (~(U2v2a4 & Wffw84));
	assign U2v2a4 = (Yq13a4 & Fr13a4);
	assign Yq13a4 = (~(Yvb2a4 | Km63a4[0]));
	assign Pp13a4 = (Mr13a4 & Tr13a4);
	assign Tr13a4 = (~(B3v2a4 & Etdw84));
	assign B3v2a4 = (As13a4 & Fr13a4);
	assign As13a4 = (~(V2vx84 | Yvb2a4));
	assign Mr13a4 = (~(K4v2a4 & Gpiw84));
	assign K4v2a4 = (Fr13a4 & Rq13a4);
	assign Bp13a4 = (~(Hs13a4 | I4g2a4));
	assign Hs13a4 = (~(Os13a4 & Vs13a4));
	assign Vs13a4 = (~(R4v2a4 & O2hw84));
	assign R4v2a4 = (Fr13a4 & Zh03a4);
	assign Fr13a4 = (~(N5vx84 | Km63a4[2]));
	assign Os13a4 = (~(F5v2a4 & Ujaw84));
	assign Tyu2a4 = (Ct13a4 & Jt13a4);
	assign Go13a4 = (~(M5v2a4 & Cx8w84));
	assign M5v2a4 = (~(M7ix84 | Ct13a4));
	assign Ct13a4 = (Qt13a4 & Xt13a4);
	assign Xt13a4 = (Eu13a4 & Lu13a4);
	assign Lu13a4 = (~(Ffox84 | G0c2a4));
	assign Ffox84 = (F2gx84 & J13x84);
	assign Eu13a4 = (B1c2a4 & Yrix84);
	assign Yrix84 = (!E3ix84);
	assign E3ix84 = (E3wx84 & Ns2x84);
	assign E3wx84 = (~(Jnix84 | Pqbx84));
	assign Jnix84 = (!Undx84);
	assign B1c2a4 = (Bqwx84 | Gz4w84);
	assign Bqwx84 = (!Ub82a4);
	assign Ub82a4 = (~(Tsix84 | Zo2x84));
	assign Qt13a4 = (Su13a4 & Zu13a4);
	assign Zu13a4 = (~(Km63a4[0] & F5v2a4));
	assign F5v2a4 = (Km63a4[1] & Gi03a4);
	assign Gi03a4 = (~(N5vx84 | Bzux84));
	assign N5vx84 = (!Km63a4[3]);
	assign Su13a4 = (Gv13a4 & Nv13a4);
	assign Nv13a4 = (Uy1y84 | Evix84);
	assign Evix84 = (!Zgxx84);
	assign Uy1y84 = (!A2ox84);
	assign A2ox84 = (Pz2x84 & Ewax84);
	assign Gv13a4 = (J9bx84 | S1dx84);
	assign S1dx84 = (!Ap52a4);
	assign Ap52a4 = (Tq2x84 & Ns2x84);
	assign J9bx84 = (!Qvax84);
	assign Qvax84 = (Fn2x84 & J13x84);
	assign Kxu2a4 = (~(Uv13a4 & Dkix84));
	assign Uv13a4 = (~(Bw13a4 & Iw13a4));
	assign Iw13a4 = (~(Pw13a4 & Ambx84));
	assign Pw13a4 = (~(Ww13a4 & Dx13a4));
	assign Dx13a4 = (Kx13a4 & Rx13a4);
	assign Rx13a4 = (~(Yx13a4 & S3ix84));
	assign Yx13a4 = (~(H8px84 | Ewax84));
	assign H8px84 = (!Drbx84);
	assign Drbx84 = (Pz2x84 & Mmvx84);
	assign Kx13a4 = (~(Jsrx84 | Q0yx84));
	assign Jsrx84 = (Y6bx84 & Bw2x84);
	assign Ww13a4 = (Fy13a4 & My13a4);
	assign My13a4 = (W1c2a4 | Yqcx84);
	assign W1c2a4 = (!Hghx84);
	assign Hghx84 = (Hu2x84 & G4bx84);
	assign Fy13a4 = (Tswx84 | Mmvx84);
	assign Tswx84 = (!Mgnx84);
	assign Mgnx84 = (Zo2x84 & Ns2x84);
	assign Bw13a4 = (Ty13a4 & O22y84);
	assign O22y84 = (~(Az13a4 & M7ix84));
	assign M7ix84 = (!Jt13a4);
	assign Az13a4 = (D8gx84 ? Oz13a4 : Hz13a4);
	assign Ty13a4 = (~(Vz13a4 & Uwix84));
	assign Uwix84 = (Yqcx84 & Mmvx84);
	assign Vz13a4 = (~(Fn2x84 | Ns2x84));
	assign Sn13a4 = (~(Qp63a4[0] & T5v2a4));
	assign T5v2a4 = (C023a4 & Dkix84);
	assign Dkix84 = (~(J023a4 & Q023a4));
	assign Q023a4 = (X023a4 & E123a4);
	assign E123a4 = (L123a4 & S123a4);
	assign S123a4 = (~(Yzhx84 & Z123a4));
	assign Z123a4 = (Krix84 | G223a4);
	assign G223a4 = (~(H6dx84 | Yqcx84));
	assign Krix84 = (D9mx84 & Ewax84);
	assign Yzhx84 = (Wqbx84 & Tsix84);
	assign L123a4 = (Q813a4 & Pd2y84);
	assign Q813a4 = (~(N223a4 & S3ix84));
	assign S3ix84 = (Zo2x84 & Fn2x84);
	assign N223a4 = (~(Fycx84 | D4dx84));
	assign Fycx84 = (!F352a4);
	assign F352a4 = (Vx2x84 & Mmvx84);
	assign X023a4 = (U223a4 & B323a4);
	assign B323a4 = (~(Gcvx84 & I323a4));
	assign I323a4 = (~(Gzfx84 & P323a4));
	assign P323a4 = (~(W323a4 & Uacx84));
	assign W323a4 = (~(Ambx84 | N4ix84));
	assign Gzfx84 = (!Q0yx84);
	assign Q0yx84 = (Hu2x84 & Bw2x84);
	assign U223a4 = (~(Tq2x84 & D423a4));
	assign D423a4 = (E1dx84 | K423a4);
	assign K423a4 = (Nacx84 & D9mx84);
	assign D9mx84 = (~(N4ix84 | J13x84));
	assign E1dx84 = (Mlbx84 & Pqbx84);
	assign J023a4 = (R423a4 & Y423a4);
	assign Y423a4 = (F523a4 & M523a4);
	assign M523a4 = (Y1d2a4 | Pqbx84);
	assign Pqbx84 = (!Pz2x84);
	assign Y1d2a4 = (~(T523a4 & Gwix84));
	assign T523a4 = (~(Zo2x84 | Ns2x84));
	assign F523a4 = (~(A623a4 & H6dx84));
	assign H6dx84 = (!D53x84);
	assign A623a4 = (~(H623a4 & O623a4));
	assign O623a4 = (~(Rzhx84 & Uacx84));
	assign Uacx84 = (~(Wqbx84 | Tq2x84));
	assign Rzhx84 = (~(Ucox84 | Vx2x84));
	assign Ucox84 = (!Phdx84);
	assign Phdx84 = (~(Fmvx84 | N4ix84));
	assign H623a4 = (V623a4 & C723a4);
	assign C723a4 = (~(J723a4 & Y1gx84));
	assign Y1gx84 = (~(Fmvx84 | D4dx84));
	assign Fmvx84 = (!Pxbx84);
	assign Pxbx84 = (Gpbx84 & Ambx84);
	assign J723a4 = (~(Yqcx84 | N4ix84));
	assign V623a4 = (~(Q723a4 & Mlbx84));
	assign Mlbx84 = (Hgvx84 & Gpbx84);
	assign Hgvx84 = (!N4ix84);
	assign Q723a4 = (Y3i2a4 & Qxmx84);
	assign R423a4 = (Uvu2a4 & E8a2a4);
	assign E8a2a4 = (X723a4 & E823a4);
	assign E823a4 = (~(L823a4 & Livx84));
	assign Livx84 = (G4bx84 & Tsix84);
	assign L823a4 = (~(B5bx84 | Gz4w84));
	assign B5bx84 = (!Sbvx84);
	assign Sbvx84 = (Hu2x84 & Vx2x84);
	assign X723a4 = (~(T613a4 & B9lx84));
	assign T613a4 = (Y3i2a4 & Undx84);
	assign Undx84 = (Mmvx84 & Qxmx84);
	assign Y3i2a4 = (~(G4bx84 | Ns2x84));
	assign Uvu2a4 = (S823a4 & Z823a4);
	assign Z823a4 = (G923a4 & N923a4);
	assign N923a4 = (~(U923a4 & Ozcx84));
	assign Ozcx84 = (Y6bx84 & Qxmx84);
	assign Y6bx84 = (Zo2x84 & Wqbx84);
	assign U923a4 = (~(Ambx84 | D53x84));
	assign Ambx84 = (!J13x84);
	assign G923a4 = (Iu42a4 & Gqox84);
	assign Gqox84 = (Fthx84 | Pz2x84);
	assign Fthx84 = (!Gcvx84);
	assign Iu42a4 = (O2ox84 | Uj2x84);
	assign O2ox84 = (~(Ba23a4 & Gwix84));
	assign Ba23a4 = (~(D4dx84 | Zo2x84));
	assign S823a4 = (Ia23a4 & Pa23a4);
	assign Pa23a4 = (Vzcx84 | Nbix84);
	assign Nbix84 = (!Wdox84);
	assign Wdox84 = (Nwix84 & Gcvx84);
	assign Nwix84 = (~(Jxmx84 | Wqbx84));
	assign Jxmx84 = (!Gwix84);
	assign Gwix84 = (J13x84 & G4bx84);
	assign Vzcx84 = (~(Wa23a4 & Db23a4));
	assign Db23a4 = (Kb23a4 & Rb23a4);
	assign Rb23a4 = (Yb23a4 & Fc23a4);
	assign Fc23a4 = (~(Xw6w84 & Mc23a4));
	assign Mc23a4 = (Iv6w84 | My6w84);
	assign Yb23a4 = (~(Pq6w84 & Tkcx84));
	assign Kb23a4 = (Tc23a4 & Ad23a4);
	assign Ad23a4 = (~(Tt6w84 & Sgcx84));
	assign Sgcx84 = (Kjcx84 | Es6w84);
	assign Tc23a4 = (~(Es6w84 & Kjcx84));
	assign Kjcx84 = (Tkcx84 | Pq6w84);
	assign Tkcx84 = (!Nlmx84);
	assign Nlmx84 = (Njox84 & D8gx84);
	assign Wa23a4 = (Hd23a4 & Od23a4);
	assign Od23a4 = (Dnmx84 | Tmox84);
	assign Dnmx84 = (!Iv6w84);
	assign Hd23a4 = (Vd23a4 & Ce23a4);
	assign Ce23a4 = (D8gx84 | Njox84);
	assign Njox84 = (Gjox84 & T7px84);
	assign D8gx84 = (!Ap6w84);
	assign Vd23a4 = (T7px84 | Gjox84);
	assign Gjox84 = (!Vfbx84);
	assign Vfbx84 = (~(Xhox84 & Tmox84));
	assign Tmox84 = (!My6w84);
	assign Xhox84 = (~(Iv6w84 | Xw6w84));
	assign T7px84 = (!C07w84);
	assign Ia23a4 = (~(Iqbx84 & Wlnx84));
	assign Wlnx84 = (Tq2x84 & Tsix84);
	assign Iqbx84 = (Gcvx84 & Qxmx84);
	assign Gcvx84 = (Zo2x84 & Ewax84);
	assign Ewax84 = (!Vx2x84);
	assign C023a4 = (~(Je23a4 & Qe23a4));
	assign Qe23a4 = (Xe23a4 & Ef23a4);
	assign Ef23a4 = (~(G0c2a4 | Lw72a4));
	assign Lw72a4 = (Tq2x84 & Wqbx84);
	assign Wqbx84 = (!Ns2x84);
	assign G0c2a4 = (Zgxx84 & Qxmx84);
	assign Zgxx84 = (Bw2x84 & Ns2x84);
	assign Xe23a4 = (~(Aq42a4 | Gc72a4));
	assign Gc72a4 = (Zo2x84 & J13x84);
	assign Aq42a4 = (Gpix84 & Zo2x84);
	assign Gpix84 = (~(Fn2x84 | Hu2x84));
	assign Je23a4 = (Lf23a4 & Sf23a4);
	assign Sf23a4 = (Zf23a4 & Iz1y84);
	assign Iz1y84 = (Gg23a4 | Jt13a4);
	assign Jt13a4 = (P7d2a4 & Ng23a4);
	assign Ng23a4 = (~(Jfxx84 & M0px84));
	assign M0px84 = (Fn2x84 & Qxmx84);
	assign Qxmx84 = (!Hu2x84);
	assign Jfxx84 = (~(Gpbx84 | D4dx84));
	assign D4dx84 = (!Xm92a4);
	assign Xm92a4 = (Ns2x84 & Tsix84);
	assign P7d2a4 = (Pd2y84 | N4ix84);
	assign N4ix84 = (Ju4w84 & Lmdx84);
	assign Lmdx84 = (!Qq8x84);
	assign Pd2y84 = (Ao62a4 | Pz2x84);
	assign Ao62a4 = (B0gx84 | Tq2x84);
	assign B0gx84 = (!B9lx84);
	assign B9lx84 = (On72a4 & Gpbx84);
	assign Gpbx84 = (!Gz4w84);
	assign On72a4 = (Vx2x84 & Yqcx84);
	assign Gg23a4 = (Ap6w84 ? Hz13a4 : Oz13a4);
	assign Hz13a4 = (Ln6w84 ? Bh23a4 : Ug23a4);
	assign Bh23a4 = (Ih23a4 & Ph23a4);
	assign Ph23a4 = (~(I3dx84 & Evf2a4));
	assign Evf2a4 = (~(Wh23a4 & Di23a4));
	assign Di23a4 = (Ki23a4 & Ri23a4);
	assign Ri23a4 = (Yi23a4 & Fj23a4);
	assign Fj23a4 = (~(Mj23a4 & Psvw84));
	assign Yi23a4 = (~(Tj23a4 & Fjsw84));
	assign Ki23a4 = (Ak23a4 & Hk23a4);
	assign Hk23a4 = (~(Ok23a4 & V9pw84));
	assign Ak23a4 = (~(Vk23a4 & L0mw84));
	assign Wh23a4 = (Cl23a4 & Jl23a4);
	assign Jl23a4 = (Ql23a4 & Xl23a4);
	assign Xl23a4 = (~(Em23a4 & X5uw84));
	assign Ql23a4 = (~(Lm23a4 & Nwqw84));
	assign Cl23a4 = (Sm23a4 & Zm23a4);
	assign Zm23a4 = (~(Gn23a4 & Dnnw84));
	assign Sm23a4 = (~(Nn23a4 & Tdkw84));
	assign Ih23a4 = (Wl6w84 ? Bo23a4 : Un23a4);
	assign Bo23a4 = (Io23a4 & Po23a4);
	assign Po23a4 = (~(Tgk2a4 & Otf2a4));
	assign Otf2a4 = (~(Wo23a4 & Dp23a4));
	assign Dp23a4 = (Kp23a4 & Rp23a4);
	assign Rp23a4 = (Yp23a4 & Fq23a4);
	assign Fq23a4 = (~(Ayvw84 & Mj23a4));
	assign Yp23a4 = (~(Qosw84 & Tj23a4));
	assign Kp23a4 = (Mq23a4 & Tq23a4);
	assign Tq23a4 = (~(Gfpw84 & Ok23a4));
	assign Mq23a4 = (~(W5mw84 & Vk23a4));
	assign Wo23a4 = (Ar23a4 & Hr23a4);
	assign Hr23a4 = (Or23a4 & Vr23a4);
	assign Vr23a4 = (~(Ibuw84 & Em23a4));
	assign Or23a4 = (~(Y1rw84 & Lm23a4));
	assign Ar23a4 = (Cs23a4 & Js23a4);
	assign Js23a4 = (~(Osnw84 & Gn23a4));
	assign Cs23a4 = (~(Ejkw84 & Nn23a4));
	assign Io23a4 = (Qs23a4 & Xs23a4);
	assign Xs23a4 = (~(Aanx84 & Vtf2a4));
	assign Vtf2a4 = (~(Et23a4 & Lt23a4));
	assign Lt23a4 = (St23a4 & Zt23a4);
	assign Zt23a4 = (Gu23a4 & Nu23a4);
	assign Nu23a4 = (~(Kuvw84 & Mj23a4));
	assign Gu23a4 = (~(Alsw84 & Tj23a4));
	assign St23a4 = (Uu23a4 & Bv23a4);
	assign Bv23a4 = (~(Qbpw84 & Ok23a4));
	assign Uu23a4 = (~(G2mw84 & Vk23a4));
	assign Et23a4 = (Iv23a4 & Pv23a4);
	assign Pv23a4 = (Wv23a4 & Dw23a4);
	assign Dw23a4 = (~(S7uw84 & Em23a4));
	assign Wv23a4 = (~(Iyqw84 & Lm23a4));
	assign Iv23a4 = (Kw23a4 & Rw23a4);
	assign Rw23a4 = (~(Yonw84 & Gn23a4));
	assign Kw23a4 = (~(Ofkw84 & Nn23a4));
	assign Qs23a4 = (~(M8ox84 & Xuf2a4));
	assign Xuf2a4 = (~(Yw23a4 & Fx23a4));
	assign Fx23a4 = (Mx23a4 & Tx23a4);
	assign Tx23a4 = (Ay23a4 & Hy23a4);
	assign Hy23a4 = (~(Fwvw84 & Mj23a4));
	assign Ay23a4 = (~(Vmsw84 & Tj23a4));
	assign Mx23a4 = (Oy23a4 & Vy23a4);
	assign Vy23a4 = (~(Ldpw84 & Ok23a4));
	assign Oy23a4 = (~(B4mw84 & Vk23a4));
	assign Yw23a4 = (Cz23a4 & Jz23a4);
	assign Jz23a4 = (Qz23a4 & Xz23a4);
	assign Xz23a4 = (~(N9uw84 & Em23a4));
	assign Qz23a4 = (~(D0rw84 & Lm23a4));
	assign Cz23a4 = (E033a4 & L033a4);
	assign L033a4 = (~(Tqnw84 & Gn23a4));
	assign E033a4 = (~(Jhkw84 & Nn23a4));
	assign Un23a4 = (S033a4 & Z033a4);
	assign Z033a4 = (G133a4 & N133a4);
	assign N133a4 = (~(Aanx84 & Ixf2a4));
	assign Ixf2a4 = (~(U133a4 & B233a4));
	assign B233a4 = (I233a4 & P233a4);
	assign P233a4 = (W233a4 & D333a4);
	assign D333a4 = (~(Q1ww84 & Mj23a4));
	assign W233a4 = (~(Gssw84 & Tj23a4));
	assign I233a4 = (K333a4 & R333a4);
	assign R333a4 = (~(Wipw84 & Ok23a4));
	assign K333a4 = (~(M9mw84 & Vk23a4));
	assign U133a4 = (Y333a4 & F433a4);
	assign F433a4 = (M433a4 & T433a4);
	assign T433a4 = (~(Yeuw84 & Em23a4));
	assign M433a4 = (~(O5rw84 & Lm23a4));
	assign Y333a4 = (A533a4 & H533a4);
	assign H533a4 = (~(Ewnw84 & Gn23a4));
	assign A533a4 = (~(Umkw84 & Nn23a4));
	assign G133a4 = (~(I0nx84 & Kyf2a4));
	assign Kyf2a4 = (~(O533a4 & V533a4));
	assign V533a4 = (C633a4 & J633a4);
	assign J633a4 = (Q633a4 & X633a4);
	assign X633a4 = (~(Vzvw84 & Mj23a4));
	assign Q633a4 = (~(Lqsw84 & Tj23a4));
	assign C633a4 = (E733a4 & L733a4);
	assign L733a4 = (~(Bhpw84 & Ok23a4));
	assign E733a4 = (~(R7mw84 & Vk23a4));
	assign O533a4 = (S733a4 & Z733a4);
	assign Z733a4 = (G833a4 & N833a4);
	assign N833a4 = (~(Dduw84 & Em23a4));
	assign G833a4 = (~(T3rw84 & Lm23a4));
	assign S733a4 = (U833a4 & B933a4);
	assign B933a4 = (~(Junw84 & Gn23a4));
	assign U833a4 = (~(Zkkw84 & Nn23a4));
	assign S033a4 = (I933a4 & P933a4);
	assign P933a4 = (~(M8ox84 & Dyf2a4));
	assign Dyf2a4 = (~(W933a4 & Da33a4));
	assign Da33a4 = (Ka33a4 & Ra33a4);
	assign Ra33a4 = (Ya33a4 & Fb33a4);
	assign Fb33a4 = (~(Mj23a4 & L3ww84));
	assign Ya33a4 = (~(Tj23a4 & Busw84));
	assign Ka33a4 = (Mb33a4 & Tb33a4);
	assign Tb33a4 = (~(Ok23a4 & Rkpw84));
	assign Mb33a4 = (~(Vk23a4 & Hbmw84));
	assign W933a4 = (Ac33a4 & Hc33a4);
	assign Hc33a4 = (Oc33a4 & Vc33a4);
	assign Vc33a4 = (~(Em23a4 & Tguw84));
	assign Oc33a4 = (~(Lm23a4 & J7rw84));
	assign Ac33a4 = (Cd33a4 & Jd33a4);
	assign Jd33a4 = (~(Gn23a4 & Zxnw84));
	assign Cd33a4 = (~(Nn23a4 & Pokw84));
	assign I933a4 = (~(Tgk2a4 & Bxf2a4));
	assign Bxf2a4 = (~(Qd33a4 & Xd33a4));
	assign Xd33a4 = (Ee33a4 & Le33a4);
	assign Le33a4 = (Se33a4 & Ze33a4);
	assign Ze33a4 = (~(G5ww84 & Mj23a4));
	assign Se33a4 = (~(Wvsw84 & Tj23a4));
	assign Ee33a4 = (Gf33a4 & Nf33a4);
	assign Nf33a4 = (~(Mmpw84 & Ok23a4));
	assign Gf33a4 = (~(Cdmw84 & Vk23a4));
	assign Qd33a4 = (Uf33a4 & Bg33a4);
	assign Bg33a4 = (Ig33a4 & Pg33a4);
	assign Pg33a4 = (~(Oiuw84 & Em23a4));
	assign Ig33a4 = (~(E9rw84 & Lm23a4));
	assign Uf33a4 = (Wg33a4 & Dh33a4);
	assign Dh33a4 = (~(Uznw84 & Gn23a4));
	assign Wg33a4 = (~(Kqkw84 & Nn23a4));
	assign Ug23a4 = (Kh33a4 & Rh33a4);
	assign Rh33a4 = (~(I3dx84 & Fdg2a4));
	assign Fdg2a4 = (~(Yh33a4 & Fi33a4));
	assign Fi33a4 = (Mi33a4 & Ti33a4);
	assign Ti33a4 = (Aj33a4 & Hj33a4);
	assign Hj33a4 = (~(B7ww84 & Mj23a4));
	assign Aj33a4 = (~(Rxsw84 & Tj23a4));
	assign Mi33a4 = (Oj33a4 & Vj33a4);
	assign Vj33a4 = (~(Hopw84 & Ok23a4));
	assign Oj33a4 = (~(Xemw84 & Vk23a4));
	assign Yh33a4 = (Ck33a4 & Jk33a4);
	assign Jk33a4 = (Qk33a4 & Xk33a4);
	assign Xk33a4 = (~(Jkuw84 & Em23a4));
	assign Qk33a4 = (~(Zarw84 & Lm23a4));
	assign Ck33a4 = (El33a4 & Ll33a4);
	assign Ll33a4 = (~(P1ow84 & Gn23a4));
	assign El33a4 = (~(Fskw84 & Nn23a4));
	assign Kh33a4 = (Wl6w84 ? Zl33a4 : Sl33a4);
	assign Zl33a4 = (Gm33a4 & Nm33a4);
	assign Nm33a4 = (~(Tgk2a4 & Wbg2a4));
	assign Wbg2a4 = (~(Um33a4 & Bn33a4));
	assign Bn33a4 = (In33a4 & Pn33a4);
	assign Pn33a4 = (Wn33a4 & Do33a4);
	assign Do33a4 = (~(Ocww84 & Mj23a4));
	assign Wn33a4 = (~(E3tw84 & Tj23a4));
	assign In33a4 = (Ko33a4 & Ro33a4);
	assign Ro33a4 = (~(Utpw84 & Ok23a4));
	assign Ko33a4 = (~(Kkmw84 & Vk23a4));
	assign Um33a4 = (Yo33a4 & Fp33a4);
	assign Fp33a4 = (Mp33a4 & Tp33a4);
	assign Tp33a4 = (~(Wpuw84 & Em23a4));
	assign Mp33a4 = (~(Mgrw84 & Lm23a4));
	assign Yo33a4 = (Aq33a4 & Hq33a4);
	assign Hq33a4 = (~(C7ow84 & Gn23a4));
	assign Aq33a4 = (~(Sxkw84 & Nn23a4));
	assign Gm33a4 = (Oq33a4 & Vq33a4);
	assign Vq33a4 = (~(Aanx84 & Dcg2a4));
	assign Dcg2a4 = (~(Cr33a4 & Jr33a4));
	assign Jr33a4 = (Qr33a4 & Xr33a4);
	assign Xr33a4 = (Es33a4 & Ls33a4);
	assign Ls33a4 = (~(W8ww84 & Mj23a4));
	assign Es33a4 = (~(Mzsw84 & Tj23a4));
	assign Qr33a4 = (Ss33a4 & Zs33a4);
	assign Zs33a4 = (~(Cqpw84 & Ok23a4));
	assign Ss33a4 = (~(Sgmw84 & Vk23a4));
	assign Cr33a4 = (Gt33a4 & Nt33a4);
	assign Nt33a4 = (Ut33a4 & Bu33a4);
	assign Bu33a4 = (~(Emuw84 & Em23a4));
	assign Ut33a4 = (~(Ucrw84 & Lm23a4));
	assign Gt33a4 = (Iu33a4 & Pu33a4);
	assign Pu33a4 = (~(K3ow84 & Gn23a4));
	assign Iu33a4 = (~(Aukw84 & Nn23a4));
	assign Oq33a4 = (~(M8ox84 & Ycg2a4));
	assign Ycg2a4 = (~(Wu33a4 & Dv33a4));
	assign Dv33a4 = (Kv33a4 & Rv33a4);
	assign Rv33a4 = (Yv33a4 & Fw33a4);
	assign Fw33a4 = (~(Saww84 & Mj23a4));
	assign Yv33a4 = (~(I1tw84 & Tj23a4));
	assign Kv33a4 = (Mw33a4 & Tw33a4);
	assign Tw33a4 = (~(Yrpw84 & Ok23a4));
	assign Mw33a4 = (~(Oimw84 & Vk23a4));
	assign Wu33a4 = (Ax33a4 & Hx33a4);
	assign Hx33a4 = (Ox33a4 & Vx33a4);
	assign Vx33a4 = (~(Aouw84 & Em23a4));
	assign Ox33a4 = (~(Qerw84 & Lm23a4));
	assign Ax33a4 = (Cy33a4 & Jy33a4);
	assign Jy33a4 = (~(G5ow84 & Gn23a4));
	assign Cy33a4 = (~(Wvkw84 & Nn23a4));
	assign Sl33a4 = (Qy33a4 & Xy33a4);
	assign Xy33a4 = (Ez33a4 & Lz33a4);
	assign Lz33a4 = (~(I0nx84 & Xfg2a4));
	assign Xfg2a4 = (~(Sz33a4 & Zz33a4));
	assign Zz33a4 = (G043a4 & N043a4);
	assign N043a4 = (U043a4 & B143a4);
	assign B143a4 = (~(Keww84 & Mj23a4));
	assign U043a4 = (~(A5tw84 & Tj23a4));
	assign G043a4 = (I143a4 & P143a4);
	assign P143a4 = (~(Qvpw84 & Ok23a4));
	assign I143a4 = (~(Gmmw84 & Vk23a4));
	assign Sz33a4 = (W143a4 & D243a4);
	assign D243a4 = (K243a4 & R243a4);
	assign R243a4 = (~(Sruw84 & Em23a4));
	assign K243a4 = (~(Iirw84 & Lm23a4));
	assign W143a4 = (Y243a4 & F343a4);
	assign F343a4 = (~(Y8ow84 & Gn23a4));
	assign Y243a4 = (~(Ozkw84 & Nn23a4));
	assign Ez33a4 = (~(Aanx84 & Veg2a4));
	assign Veg2a4 = (~(M343a4 & T343a4));
	assign T343a4 = (A443a4 & H443a4);
	assign H443a4 = (O443a4 & V443a4);
	assign V443a4 = (~(Ggww84 & Mj23a4));
	assign O443a4 = (~(W6tw84 & Tj23a4));
	assign A443a4 = (C543a4 & J543a4);
	assign J543a4 = (~(Mxpw84 & Ok23a4));
	assign C543a4 = (~(Comw84 & Vk23a4));
	assign M343a4 = (Q543a4 & X543a4);
	assign X543a4 = (E643a4 & L643a4);
	assign L643a4 = (~(Otuw84 & Em23a4));
	assign E643a4 = (~(Ekrw84 & Lm23a4));
	assign Q543a4 = (S643a4 & Z643a4);
	assign Z643a4 = (~(Uaow84 & Gn23a4));
	assign S643a4 = (~(K1lw84 & Nn23a4));
	assign Qy33a4 = (G743a4 & N743a4);
	assign N743a4 = (~(Tgk2a4 & Oeg2a4));
	assign Oeg2a4 = (~(U743a4 & B843a4));
	assign B843a4 = (I843a4 & P843a4);
	assign P843a4 = (W843a4 & D943a4);
	assign D943a4 = (~(Yjww84 & Mj23a4));
	assign W843a4 = (~(Oatw84 & Tj23a4));
	assign I843a4 = (K943a4 & R943a4);
	assign R943a4 = (~(E1qw84 & Ok23a4));
	assign K943a4 = (~(Urmw84 & Vk23a4));
	assign U743a4 = (Y943a4 & Fa43a4);
	assign Fa43a4 = (Ma43a4 & Ta43a4);
	assign Ta43a4 = (~(Gxuw84 & Em23a4));
	assign Ma43a4 = (~(Wnrw84 & Lm23a4));
	assign Y943a4 = (Ab43a4 & Hb43a4);
	assign Hb43a4 = (~(Meow84 & Gn23a4));
	assign Ab43a4 = (~(C5lw84 & Nn23a4));
	assign G743a4 = (~(M8ox84 & Qfg2a4));
	assign Qfg2a4 = (~(Ob43a4 & Vb43a4));
	assign Vb43a4 = (Cc43a4 & Jc43a4);
	assign Jc43a4 = (Qc43a4 & Xc43a4);
	assign Xc43a4 = (~(Mj23a4 & Ciww84));
	assign Qc43a4 = (~(Tj23a4 & S8tw84));
	assign Cc43a4 = (Ed43a4 & Ld43a4);
	assign Ld43a4 = (~(Ok23a4 & Izpw84));
	assign Ed43a4 = (~(Vk23a4 & Ypmw84));
	assign Ob43a4 = (Sd43a4 & Zd43a4);
	assign Zd43a4 = (Ge43a4 & Ne43a4);
	assign Ne43a4 = (~(Em23a4 & Kvuw84));
	assign Ge43a4 = (~(Lm23a4 & Amrw84));
	assign Sd43a4 = (Ue43a4 & Bf43a4);
	assign Bf43a4 = (~(Gn23a4 & Qcow84));
	assign Ue43a4 = (~(Nn23a4 & G3lw84));
	assign Oz13a4 = (Ln6w84 ? Pf43a4 : If43a4);
	assign Pf43a4 = (Wf43a4 & Dg43a4);
	assign Dg43a4 = (~(I3dx84 & Cmg2a4));
	assign Cmg2a4 = (~(Kg43a4 & Rg43a4));
	assign Rg43a4 = (Yg43a4 & Fh43a4);
	assign Fh43a4 = (Mh43a4 & Th43a4);
	assign Th43a4 = (~(Ulww84 & Mj23a4));
	assign Mh43a4 = (~(Kctw84 & Tj23a4));
	assign Yg43a4 = (Ai43a4 & Hi43a4);
	assign Hi43a4 = (~(A3qw84 & Ok23a4));
	assign Ai43a4 = (~(Qtmw84 & Vk23a4));
	assign Kg43a4 = (Oi43a4 & Vi43a4);
	assign Vi43a4 = (Cj43a4 & Jj43a4);
	assign Jj43a4 = (~(Czuw84 & Em23a4));
	assign Cj43a4 = (~(Sprw84 & Lm23a4));
	assign Oi43a4 = (Qj43a4 & Xj43a4);
	assign Xj43a4 = (~(Igow84 & Gn23a4));
	assign Qj43a4 = (~(Y6lw84 & Nn23a4));
	assign Wf43a4 = (Wl6w84 ? Lk43a4 : Ek43a4);
	assign Lk43a4 = (Sk43a4 & Zk43a4);
	assign Zk43a4 = (~(Tgk2a4 & Tkg2a4));
	assign Tkg2a4 = (~(Gl43a4 & Nl43a4));
	assign Nl43a4 = (Ul43a4 & Bm43a4);
	assign Bm43a4 = (Im43a4 & Pm43a4);
	assign Pm43a4 = (~(Irww84 & Mj23a4));
	assign Im43a4 = (~(Yhtw84 & Tj23a4));
	assign Ul43a4 = (Wm43a4 & Dn43a4);
	assign Dn43a4 = (~(O8qw84 & Ok23a4));
	assign Wm43a4 = (~(Ezmw84 & Vk23a4));
	assign Gl43a4 = (Kn43a4 & Rn43a4);
	assign Rn43a4 = (Yn43a4 & Fo43a4);
	assign Fo43a4 = (~(Q4vw84 & Em23a4));
	assign Yn43a4 = (~(Gvrw84 & Lm23a4));
	assign Kn43a4 = (Mo43a4 & To43a4);
	assign To43a4 = (~(Wlow84 & Gn23a4));
	assign Mo43a4 = (~(Mclw84 & Nn23a4));
	assign Sk43a4 = (Ap43a4 & Hp43a4);
	assign Hp43a4 = (~(Aanx84 & Alg2a4));
	assign Alg2a4 = (~(Op43a4 & Vp43a4));
	assign Vp43a4 = (Cq43a4 & Jq43a4);
	assign Jq43a4 = (Qq43a4 & Xq43a4);
	assign Xq43a4 = (~(Qnww84 & Mj23a4));
	assign Qq43a4 = (~(Getw84 & Tj23a4));
	assign Cq43a4 = (Er43a4 & Lr43a4);
	assign Lr43a4 = (~(W4qw84 & Ok23a4));
	assign Er43a4 = (~(Mvmw84 & Vk23a4));
	assign Op43a4 = (Sr43a4 & Zr43a4);
	assign Zr43a4 = (Gs43a4 & Ns43a4);
	assign Ns43a4 = (~(Y0vw84 & Em23a4));
	assign Gs43a4 = (~(Orrw84 & Lm23a4));
	assign Sr43a4 = (Us43a4 & Bt43a4);
	assign Bt43a4 = (~(Eiow84 & Gn23a4));
	assign Us43a4 = (~(U8lw84 & Nn23a4));
	assign Ap43a4 = (~(M8ox84 & Vlg2a4));
	assign Vlg2a4 = (~(It43a4 & Pt43a4));
	assign Pt43a4 = (Wt43a4 & Du43a4);
	assign Du43a4 = (Ku43a4 & Ru43a4);
	assign Ru43a4 = (~(Mpww84 & Mj23a4));
	assign Ku43a4 = (~(Cgtw84 & Tj23a4));
	assign Wt43a4 = (Yu43a4 & Fv43a4);
	assign Fv43a4 = (~(S6qw84 & Ok23a4));
	assign Yu43a4 = (~(Ixmw84 & Vk23a4));
	assign It43a4 = (Mv43a4 & Tv43a4);
	assign Tv43a4 = (Aw43a4 & Hw43a4);
	assign Hw43a4 = (~(U2vw84 & Em23a4));
	assign Aw43a4 = (~(Ktrw84 & Lm23a4));
	assign Mv43a4 = (Ow43a4 & Vw43a4);
	assign Vw43a4 = (~(Akow84 & Gn23a4));
	assign Ow43a4 = (~(Qalw84 & Nn23a4));
	assign Ek43a4 = (Cx43a4 & Jx43a4);
	assign Jx43a4 = (Qx43a4 & Xx43a4);
	assign Xx43a4 = (~(Aanx84 & Sng2a4));
	assign Sng2a4 = (~(Ey43a4 & Ly43a4));
	assign Ly43a4 = (Sy43a4 & Zy43a4);
	assign Zy43a4 = (Gz43a4 & Nz43a4);
	assign Nz43a4 = (~(Avww84 & Mj23a4));
	assign Gz43a4 = (~(Qltw84 & Tj23a4));
	assign Sy43a4 = (Uz43a4 & B053a4);
	assign B053a4 = (~(Gcqw84 & Ok23a4));
	assign Uz43a4 = (~(W2nw84 & Vk23a4));
	assign Ey43a4 = (I053a4 & P053a4);
	assign P053a4 = (W053a4 & D153a4);
	assign D153a4 = (~(I8vw84 & Em23a4));
	assign W053a4 = (~(Yyrw84 & Lm23a4));
	assign I053a4 = (K153a4 & R153a4);
	assign R153a4 = (~(Opow84 & Gn23a4));
	assign K153a4 = (~(Eglw84 & Nn23a4));
	assign Qx43a4 = (~(I0nx84 & Uog2a4));
	assign Uog2a4 = (~(Y153a4 & F253a4));
	assign F253a4 = (M253a4 & T253a4);
	assign T253a4 = (A353a4 & H353a4);
	assign H353a4 = (~(Etww84 & Mj23a4));
	assign A353a4 = (~(Ujtw84 & Tj23a4));
	assign M253a4 = (O353a4 & V353a4);
	assign V353a4 = (~(Kaqw84 & Ok23a4));
	assign O353a4 = (~(A1nw84 & Vk23a4));
	assign Y153a4 = (C453a4 & J453a4);
	assign J453a4 = (Q453a4 & X453a4);
	assign X453a4 = (~(M6vw84 & Em23a4));
	assign Q453a4 = (~(Cxrw84 & Lm23a4));
	assign C453a4 = (E553a4 & L553a4);
	assign L553a4 = (~(Snow84 & Gn23a4));
	assign E553a4 = (~(Ielw84 & Nn23a4));
	assign Cx43a4 = (S553a4 & Z553a4);
	assign Z553a4 = (~(Tgk2a4 & Lng2a4));
	assign Lng2a4 = (~(G653a4 & N653a4));
	assign N653a4 = (U653a4 & B753a4);
	assign B753a4 = (I753a4 & P753a4);
	assign P753a4 = (~(Syww84 & Mj23a4));
	assign I753a4 = (~(Iptw84 & Tj23a4));
	assign U653a4 = (W753a4 & D853a4);
	assign D853a4 = (~(Yfqw84 & Ok23a4));
	assign W753a4 = (~(O6nw84 & Vk23a4));
	assign G653a4 = (K853a4 & R853a4);
	assign R853a4 = (Y853a4 & F953a4);
	assign F953a4 = (~(Acvw84 & Em23a4));
	assign Y853a4 = (~(Q2sw84 & Lm23a4));
	assign K853a4 = (M953a4 & T953a4);
	assign T953a4 = (~(Gtow84 & Gn23a4));
	assign M953a4 = (~(Wjlw84 & Nn23a4));
	assign S553a4 = (~(M8ox84 & Nog2a4));
	assign Nog2a4 = (~(Aa53a4 & Ha53a4));
	assign Ha53a4 = (Oa53a4 & Va53a4);
	assign Va53a4 = (Cb53a4 & Jb53a4);
	assign Jb53a4 = (~(Wwww84 & Mj23a4));
	assign Cb53a4 = (~(Mntw84 & Tj23a4));
	assign Oa53a4 = (Qb53a4 & Xb53a4);
	assign Xb53a4 = (~(Ceqw84 & Ok23a4));
	assign Qb53a4 = (~(S4nw84 & Vk23a4));
	assign Aa53a4 = (Ec53a4 & Lc53a4);
	assign Lc53a4 = (Sc53a4 & Zc53a4);
	assign Zc53a4 = (~(Eavw84 & Em23a4));
	assign Sc53a4 = (~(U0sw84 & Lm23a4));
	assign Ec53a4 = (Gd53a4 & Nd53a4);
	assign Nd53a4 = (~(Krow84 & Gn23a4));
	assign Gd53a4 = (~(Ailw84 & Nn23a4));
	assign If43a4 = (Ud53a4 & Be53a4);
	assign Be53a4 = (~(I3dx84 & J8g2a4));
	assign J8g2a4 = (~(Ie53a4 & Pe53a4));
	assign Pe53a4 = (We53a4 & Df53a4);
	assign Df53a4 = (Kf53a4 & Rf53a4);
	assign Rf53a4 = (~(O0xw84 & Mj23a4));
	assign Kf53a4 = (~(Ertw84 & Tj23a4));
	assign We53a4 = (Yf53a4 & Fg53a4);
	assign Fg53a4 = (~(Uhqw84 & Ok23a4));
	assign Yf53a4 = (~(K8nw84 & Vk23a4));
	assign Ie53a4 = (Mg53a4 & Tg53a4);
	assign Tg53a4 = (Ah53a4 & Hh53a4);
	assign Hh53a4 = (~(Wdvw84 & Em23a4));
	assign Ah53a4 = (~(M4sw84 & Lm23a4));
	assign Mg53a4 = (Oh53a4 & Vh53a4);
	assign Vh53a4 = (~(Cvow84 & Gn23a4));
	assign Oh53a4 = (~(Sllw84 & Nn23a4));
	assign I3dx84 = (I0nx84 & Wl6w84);
	assign Ud53a4 = (Wl6w84 ? Ji53a4 : Ci53a4);
	assign Ji53a4 = (Qi53a4 & Xi53a4);
	assign Xi53a4 = (~(Tgk2a4 & A7g2a4));
	assign A7g2a4 = (~(Ej53a4 & Lj53a4));
	assign Lj53a4 = (Sj53a4 & Zj53a4);
	assign Zj53a4 = (Gk53a4 & Nk53a4);
	assign Nk53a4 = (~(C6xw84 & Mj23a4));
	assign Gk53a4 = (~(Swtw84 & Tj23a4));
	assign Sj53a4 = (Uk53a4 & Bl53a4);
	assign Bl53a4 = (~(Inqw84 & Ok23a4));
	assign Uk53a4 = (~(Ydnw84 & Vk23a4));
	assign Ej53a4 = (Il53a4 & Pl53a4);
	assign Pl53a4 = (Wl53a4 & Dm53a4);
	assign Dm53a4 = (~(Kjvw84 & Em23a4));
	assign Wl53a4 = (~(Aasw84 & Lm23a4));
	assign Il53a4 = (Km53a4 & Rm53a4);
	assign Rm53a4 = (~(Q0pw84 & Gn23a4));
	assign Km53a4 = (~(Grlw84 & Nn23a4));
	assign Qi53a4 = (Ym53a4 & Fn53a4);
	assign Fn53a4 = (~(Aanx84 & H7g2a4));
	assign H7g2a4 = (~(Mn53a4 & Tn53a4));
	assign Tn53a4 = (Ao53a4 & Ho53a4);
	assign Ho53a4 = (Oo53a4 & Vo53a4);
	assign Vo53a4 = (~(Mj23a4 & K2xw84));
	assign Oo53a4 = (~(Tj23a4 & Attw84));
	assign Ao53a4 = (Cp53a4 & Jp53a4);
	assign Jp53a4 = (~(Ok23a4 & Qjqw84));
	assign Cp53a4 = (~(Vk23a4 & Ganw84));
	assign Mn53a4 = (Qp53a4 & Xp53a4);
	assign Xp53a4 = (Eq53a4 & Lq53a4);
	assign Lq53a4 = (~(Em23a4 & Sfvw84));
	assign Eq53a4 = (~(Lm23a4 & I6sw84));
	assign Qp53a4 = (Sq53a4 & Zq53a4);
	assign Zq53a4 = (~(Gn23a4 & Ywow84));
	assign Sq53a4 = (~(Nn23a4 & Onlw84));
	assign Ym53a4 = (~(M8ox84 & C8g2a4));
	assign C8g2a4 = (~(Gr53a4 & Nr53a4));
	assign Nr53a4 = (Ur53a4 & Bs53a4);
	assign Bs53a4 = (Is53a4 & Ps53a4);
	assign Ps53a4 = (~(G4xw84 & Mj23a4));
	assign Is53a4 = (~(Wutw84 & Tj23a4));
	assign Ur53a4 = (Ws53a4 & Dt53a4);
	assign Dt53a4 = (~(Mlqw84 & Ok23a4));
	assign Ws53a4 = (~(Ccnw84 & Vk23a4));
	assign Gr53a4 = (Kt53a4 & Rt53a4);
	assign Rt53a4 = (Yt53a4 & Fu53a4);
	assign Fu53a4 = (~(Ohvw84 & Em23a4));
	assign Yt53a4 = (~(E8sw84 & Lm23a4));
	assign Kt53a4 = (Mu53a4 & Tu53a4);
	assign Tu53a4 = (~(Uyow84 & Gn23a4));
	assign Mu53a4 = (~(Kplw84 & Nn23a4));
	assign Ci53a4 = (Av53a4 & Hv53a4);
	assign Hv53a4 = (Ov53a4 & Vv53a4);
	assign Vv53a4 = (~(Aanx84 & P4g2a4));
	assign P4g2a4 = (~(Cw53a4 & Jw53a4));
	assign Jw53a4 = (Qw53a4 & Xw53a4);
	assign Xw53a4 = (Ex53a4 & Lx53a4);
	assign Lx53a4 = (~(U9xw84 & Mj23a4));
	assign Ex53a4 = (~(K0uw84 & Tj23a4));
	assign Qw53a4 = (Sx53a4 & Zx53a4);
	assign Zx53a4 = (~(Arqw84 & Ok23a4));
	assign Sx53a4 = (~(Qhnw84 & Vk23a4));
	assign Cw53a4 = (Gy53a4 & Ny53a4);
	assign Ny53a4 = (Uy53a4 & Bz53a4);
	assign Bz53a4 = (~(Cnvw84 & Em23a4));
	assign Uy53a4 = (~(Sdsw84 & Lm23a4));
	assign Gy53a4 = (Iz53a4 & Pz53a4);
	assign Pz53a4 = (~(I4pw84 & Gn23a4));
	assign Iz53a4 = (~(Yulw84 & Nn23a4));
	assign Aanx84 = (~(Hanx84 | Si6w84));
	assign Hanx84 = (!Hk6w84);
	assign Ov53a4 = (~(I0nx84 & R5g2a4));
	assign R5g2a4 = (~(Wz53a4 & D063a4));
	assign D063a4 = (K063a4 & R063a4);
	assign R063a4 = (Y063a4 & F163a4);
	assign F163a4 = (~(Y7xw84 & Mj23a4));
	assign Y063a4 = (~(Oytw84 & Tj23a4));
	assign K063a4 = (M163a4 & T163a4);
	assign T163a4 = (~(Epqw84 & Ok23a4));
	assign M163a4 = (~(Ufnw84 & Vk23a4));
	assign Wz53a4 = (A263a4 & H263a4);
	assign H263a4 = (O263a4 & V263a4);
	assign V263a4 = (~(Glvw84 & Em23a4));
	assign O263a4 = (~(Wbsw84 & Lm23a4));
	assign A263a4 = (C363a4 & J363a4);
	assign J363a4 = (~(M2pw84 & Gn23a4));
	assign C363a4 = (~(Ctlw84 & Nn23a4));
	assign I0nx84 = (Si6w84 & Hk6w84);
	assign Av53a4 = (Q363a4 & X363a4);
	assign X363a4 = (~(Tgk2a4 & I4g2a4));
	assign I4g2a4 = (~(E463a4 & L463a4));
	assign L463a4 = (S463a4 & Z463a4);
	assign Z463a4 = (G563a4 & N563a4);
	assign N563a4 = (~(Mj23a4 & Uqvw84));
	assign G563a4 = (~(Tj23a4 & Khsw84));
	assign S463a4 = (U563a4 & B663a4);
	assign B663a4 = (~(Ok23a4 & A8pw84));
	assign U563a4 = (~(Vk23a4 & Qylw84));
	assign E463a4 = (I663a4 & P663a4);
	assign P663a4 = (W663a4 & D763a4);
	assign D763a4 = (~(Em23a4 & C4uw84));
	assign W663a4 = (~(Lm23a4 & Suqw84));
	assign I663a4 = (K763a4 & R763a4);
	assign R763a4 = (~(Gn23a4 & Ilnw84));
	assign K763a4 = (~(Nn23a4 & Ybkw84));
	assign Tgk2a4 = (~(Si6w84 | Hk6w84));
	assign Q363a4 = (~(M8ox84 & K5g2a4));
	assign K5g2a4 = (~(Y763a4 & F863a4));
	assign F863a4 = (M863a4 & T863a4);
	assign T863a4 = (A963a4 & H963a4);
	assign H963a4 = (~(Mj23a4 & Qbxw84));
	assign Mj23a4 = (O963a4 & Rq13a4);
	assign A963a4 = (~(Tj23a4 & G2uw84));
	assign Tj23a4 = (V963a4 & Ca63a4);
	assign V963a4 = (~(Km63a4[0] | Km63a4[2]));
	assign M863a4 = (Ja63a4 & Qa63a4);
	assign Qa63a4 = (~(Ok23a4 & Wsqw84));
	assign Ok23a4 = (Xa63a4 & Rq13a4);
	assign Rq13a4 = (~(Km63a4[0] | Km63a4[1]));
	assign Ja63a4 = (~(Vk23a4 & Mjnw84));
	assign Vk23a4 = (Eb63a4 & Ca63a4);
	assign Eb63a4 = (~(Bzux84 | Km63a4[0]));
	assign Y763a4 = (Lb63a4 & Sb63a4);
	assign Sb63a4 = (Zb63a4 & Gc63a4);
	assign Gc63a4 = (~(Em23a4 & Yovw84));
	assign Em23a4 = (O963a4 & Zh03a4);
	assign O963a4 = (~(Km63a4[2] | Km63a4[3]));
	assign Zb63a4 = (~(Lm23a4 & Ofsw84));
	assign Lm23a4 = (Nc63a4 & Ca63a4);
	assign Nc63a4 = (~(V2vx84 | Km63a4[2]));
	assign Lb63a4 = (Uc63a4 & Bd63a4);
	assign Bd63a4 = (~(Gn23a4 & E6pw84));
	assign Gn23a4 = (Xa63a4 & Zh03a4);
	assign Zh03a4 = (~(V2vx84 | Km63a4[1]));
	assign Xa63a4 = (~(Bzux84 | Km63a4[3]));
	assign Uc63a4 = (~(Nn23a4 & Uwlw84));
	assign Nn23a4 = (Id63a4 & Ca63a4);
	assign Ca63a4 = (~(Yvb2a4 | Km63a4[3]));
	assign Yvb2a4 = (!Km63a4[1]);
	assign Id63a4 = (~(V2vx84 | Bzux84));
	assign Bzux84 = (!Km63a4[2]);
	assign V2vx84 = (!Km63a4[0]);
	assign M8ox84 = (~(Tn1y84 | Hk6w84));
	assign Tn1y84 = (!Si6w84);
	assign Zf23a4 = (~(Pd63a4 & Bdox84));
	assign Bdox84 = (!Kprx84);
	assign Kprx84 = (Fn2x84 & Ns2x84);
	assign Pd63a4 = (F2gx84 | Deox84);
	assign Deox84 = (Ns2x84 & Yqcx84);
	assign F2gx84 = (Fn2x84 & Yqcx84);
	assign Lf23a4 = (Wd63a4 & De63a4);
	assign De63a4 = (~(Nacx84 & Tsix84));
	assign Tsix84 = (!Bw2x84);
	assign Nacx84 = (~(G4bx84 | Vx2x84));
	assign G4bx84 = (!Fn2x84);
	assign Wd63a4 = (Yqcx84 ? Mmvx84 : Pz2x84);
	assign Yqcx84 = (!Zo2x84);
	assign Mmvx84 = (!Tq2x84);

	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Db73a4 <= 1'b0;
	end
	else
	  begin
	    Db73a4 <= Kk8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ed73a4 <= 1'b1;
	end
	else
	  begin
	    Ed73a4 <= Cr8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cf73a4 <= 1'b1;
	end
	else
	  begin
	    Cf73a4 <= Gm8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Bh73a4 <= 1'b0;
	end
	else
	  begin
	    Bh73a4 <= M18x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Aj73a4 <= 1'b0;
	end
	else
	  begin
	    Aj73a4 <= Kn8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Yk73a4 <= 1'b0;
	end
	else
	  begin
	    Yk73a4 <= Wq8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Um73a4 <= 1'b1;
	end
	else
	  begin
	    Um73a4 <= Of4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xo73a4 <= 1'b1;
	end
	else
	  begin
	    Xo73a4 <= Et7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Wq73a4 <= 1'b1;
	end
	else
	  begin
	    Wq73a4 <= Eh4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ws73a4 <= 1'b1;
	end
	else
	  begin
	    Ws73a4 <= Sp8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Qu73a4 <= 1'b1;
	end
	else
	  begin
	    Qu73a4 <= If4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Lw73a4 <= 1'b0;
	end
	else
	  begin
	    Lw73a4 <= Ms4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Fy73a4 <= 1'b1;
	end
	else
	  begin
	    Fy73a4 <= Gs4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  F083a4 <= 1'b1;
	end
	else
	  begin
	    F083a4 <= Mp4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  F283a4 <= 1'b1;
	end
	else
	  begin
	    F283a4 <= Uo4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  F483a4 <= 1'b0;
	end
	else
	  begin
	    F483a4 <= Ebax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  B683a4 <= 1'b1;
	end
	else
	  begin
	    B683a4 <= Yv6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  A883a4 <= 1'b1;
	end
	else
	  begin
	    A883a4 <= Et6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Z983a4 <= 1'b1;
	end
	else
	  begin
	    Z983a4 <= Gs6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Yb83a4 <= 1'b1;
	end
	else
	  begin
	    Yb83a4 <= Gy7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Vd83a4 <= 1'b1;
	end
	else
	  begin
	    Vd83a4 <= Njax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Vf83a4 <= 1'b1;
	end
	else
	  begin
	    Vf83a4 <= M15x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Vh83a4 <= 1'b1;
	end
	else
	  begin
	    Vh83a4 <= A15x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Vj83a4 <= 1'b1;
	end
	else
	  begin
	    Vj83a4 <= Qt4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Vl83a4 <= 1'b1;
	end
	else
	  begin
	    Vl83a4 <= Ys4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Vn83a4 <= 1'b0;
	end
	else
	  begin
	    Vn83a4 <= W58x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Sp83a4 <= 1'b1;
	end
	else
	  begin
	    Sp83a4 <= Xoax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rr83a4 <= 1'b1;
	end
	else
	  begin
	    Rr83a4 <= Zbax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Nt83a4 <= 1'b0;
	end
	else
	  begin
	    Nt83a4 <= A18x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Kv83a4 <= 1'b0;
	end
	else
	  begin
	    Kv83a4 <= Yi3x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hx83a4 <= 1'b1;
	end
	else
	  begin
	    Hx83a4 <= Epax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Gz83a4 <= 1'b1;
	end
	else
	  begin
	    Gz83a4 <= Cu7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  F193a4 <= 1'b1;
	end
	else
	  begin
	    F193a4 <= Gs8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  I393a4 <= 1'b1;
	end
	else
	  begin
	    I393a4 <= Lpax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  H593a4 <= 1'b1;
	end
	else
	  begin
	    H593a4 <= Iu7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  G793a4 <= 1'b0;
	end
	else
	  begin
	    G793a4 <= Cf4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  E993a4 <= 1'b0;
	end
	else
	  begin
	    E993a4 <= We4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cb93a4 <= 1'b0;
	end
	else
	  begin
	    Cb93a4 <= Qe4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ad93a4 <= 1'b1;
	end
	else
	  begin
	    Ad93a4 <= Ke4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ve93a4 <= 1'b1;
	end
	else
	  begin
	    Ve93a4 <= Q58x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rg93a4 <= 1'b1;
	end
	else
	  begin
	    Rg93a4 <= M17x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Qi93a4 <= 1'b1;
	end
	else
	  begin
	    Qi93a4 <= Q27x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Pk93a4 <= 1'b1;
	end
	else
	  begin
	    Pk93a4 <= S17x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Om93a4 <= 1'b1;
	end
	else
	  begin
	    Om93a4 <= Eq8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Lo93a4 <= 1'b1;
	end
	else
	  begin
	    Lo93a4 <= En8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Lq93a4 <= 1'b0;
	end
	else
	  begin
	    Lq93a4 <= E88x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ms93a4 <= 1'b1;
	end
	else
	  begin
	    Ms93a4 <= Ee4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mu93a4 <= 1'b1;
	end
	else
	  begin
	    Mu93a4 <= Av7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Nw93a4 <= 1'b0;
	end
	else
	  begin
	    Nw93a4 <= Yd4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ly93a4 <= 1'b0;
	end
	else
	  begin
	    Ly93a4 <= As8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  J0a3a4 <= 1'b0;
	end
	else
	  begin
	    J0a3a4 <= Sd4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  H2a3a4 <= 1'b0;
	end
	else
	  begin
	    H2a3a4 <= Il8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  D4a3a4 <= 1'b1;
	end
	else
	  begin
	    D4a3a4 <= Mm8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Z5a3a4 <= 1'b1;
	end
	else
	  begin
	    Z5a3a4 <= Ee8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  B8a3a4 <= 1'b1;
	end
	else
	  begin
	    B8a3a4 <= Mfax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Daa3a4 <= 1'b1;
	end
	else
	  begin
	    Daa3a4 <= Aa7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cca3a4 <= 1'b1;
	end
	else
	  begin
	    Cca3a4 <= Cl8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Bea3a4 <= 1'b1;
	end
	else
	  begin
	    Bea3a4 <= Co4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Yfa3a4 <= 1'b1;
	end
	else
	  begin
	    Yfa3a4 <= Ylax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Yha3a4 <= 1'b1;
	end
	else
	  begin
	    Yha3a4 <= Of8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Aka3a4 <= 1'b1;
	end
	else
	  begin
	    Aka3a4 <= Chax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cma3a4 <= 1'b0;
	end
	else
	  begin
	    Cma3a4 <= S78x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Boa3a4 <= 1'b1;
	end
	else
	  begin
	    Boa3a4 <= Gp8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Upa3a4 <= 1'b1;
	end
	else
	  begin
	    Upa3a4 <= Qoax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Tra3a4 <= 1'b0;
	end
	else
	  begin
	    Tra3a4 <= G78x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Pta3a4 <= 1'b1;
	end
	else
	  begin
	    Pta3a4 <= Ur6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mva3a4 <= 1'b1;
	end
	else
	  begin
	    Mva3a4 <= Wkax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mxa3a4 <= 1'b1;
	end
	else
	  begin
	    Mxa3a4 <= Mg8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Oza3a4 <= 1'b1;
	end
	else
	  begin
	    Oza3a4 <= Eiax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Q1b3a4 <= 1'b1;
	end
	else
	  begin
	    Q1b3a4 <= As6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  N3b3a4 <= 1'b1;
	end
	else
	  begin
	    N3b3a4 <= Anax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  N5b3a4 <= 1'b1;
	end
	else
	  begin
	    N5b3a4 <= Qe8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  P7b3a4 <= 1'b1;
	end
	else
	  begin
	    P7b3a4 <= Agax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  R9b3a4 <= 1'b1;
	end
	else
	  begin
	    R9b3a4 <= Mg5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rbb3a4 <= 1'b1;
	end
	else
	  begin
	    Rbb3a4 <= Ag5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rdb3a4 <= 1'b1;
	end
	else
	  begin
	    Rdb3a4 <= Uf4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Lfb3a4 <= 1'b1;
	end
	else
	  begin
	    Lfb3a4 <= I97x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Lhb3a4 <= 1'b1;
	end
	else
	  begin
	    Lhb3a4 <= Io4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ljb3a4 <= 1'b1;
	end
	else
	  begin
	    Ljb3a4 <= A78x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ilb3a4 <= 1'b1;
	end
	else
	  begin
	    Ilb3a4 <= Md4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Dnb3a4 <= 1'b1;
	end
	else
	  begin
	    Dnb3a4 <= Y48x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cpb3a4 <= 1'b1;
	end
	else
	  begin
	    Cpb3a4 <= Gv5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Crb3a4 <= 1'b1;
	end
	else
	  begin
	    Crb3a4 <= Uu5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ctb3a4 <= 1'b0;
	end
	else
	  begin
	    Ctb3a4 <= Ya8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Dvb3a4 <= 1'b1;
	end
	else
	  begin
	    Dvb3a4 <= G48x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Axb3a4 <= 1'b1;
	end
	else
	  begin
	    Axb3a4 <= Fmax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Azb3a4 <= 1'b1;
	end
	else
	  begin
	    Azb3a4 <= Il4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  A1c3a4 <= 1'b1;
	end
	else
	  begin
	    A1c3a4 <= Qk4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  A3c3a4 <= 1'b1;
	end
	else
	  begin
	    A3c3a4 <= G17x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  X4c3a4 <= 1'b1;
	end
	else
	  begin
	    X4c3a4 <= Hnax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  X6c3a4 <= 1'b1;
	end
	else
	  begin
	    X6c3a4 <= Ke8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Z8c3a4 <= 1'b1;
	end
	else
	  begin
	    Z8c3a4 <= Tfax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Bbc3a4 <= 1'b1;
	end
	else
	  begin
	    Bbc3a4 <= Ziax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ddc3a4 <= 1'b1;
	end
	else
	  begin
	    Ddc3a4 <= Uo6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cfc3a4 <= 1'b1;
	end
	else
	  begin
	    Cfc3a4 <= C68x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Bhc3a4 <= 1'b0;
	end
	else
	  begin
	    Bhc3a4 <= Kb8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cjc3a4 <= 1'b1;
	end
	else
	  begin
	    Cjc3a4 <= Spax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Blc3a4 <= 1'b1;
	end
	else
	  begin
	    Blc3a4 <= Uu7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Anc3a4 <= 1'b0;
	end
	else
	  begin
	    Anc3a4 <= Gd4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Yoc3a4 <= 1'b1;
	end
	else
	  begin
	    Yoc3a4 <= Ms8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Brc3a4 <= 1'b1;
	end
	else
	  begin
	    Brc3a4 <= As7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Atc3a4 <= 1'b1;
	end
	else
	  begin
	    Atc3a4 <= My7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xuc3a4 <= 1'b1;
	end
	else
	  begin
	    Xuc3a4 <= Klax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xwc3a4 <= 1'b1;
	end
	else
	  begin
	    Xwc3a4 <= Ag8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Zyc3a4 <= 1'b1;
	end
	else
	  begin
	    Zyc3a4 <= Qhax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  B1d3a4 <= 1'b1;
	end
	else
	  begin
	    B1d3a4 <= Sy7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  X2d3a4 <= 1'b1;
	end
	else
	  begin
	    X2d3a4 <= Onax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  X4d3a4 <= 1'b1;
	end
	else
	  begin
	    X4d3a4 <= Sd6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  X6d3a4 <= 1'b1;
	end
	else
	  begin
	    X6d3a4 <= Gd6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  X8d3a4 <= 1'b0;
	end
	else
	  begin
	    X8d3a4 <= Wn8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Yad3a4 <= 1'b1;
	end
	else
	  begin
	    Yad3a4 <= Ga7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xcd3a4 <= 1'b1;
	end
	else
	  begin
	    Xcd3a4 <= Uf8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Zed3a4 <= 1'b1;
	end
	else
	  begin
	    Zed3a4 <= Jhax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Bhd3a4 <= 1'b1;
	end
	else
	  begin
	    Bhd3a4 <= I08x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Yid3a4 <= 1'b1;
	end
	else
	  begin
	    Yid3a4 <= Rlax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ykd3a4 <= 1'b1;
	end
	else
	  begin
	    Ykd3a4 <= Or5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ymd3a4 <= 1'b1;
	end
	else
	  begin
	    Ymd3a4 <= Wq5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Yod3a4 <= 1'b1;
	end
	else
	  begin
	    Yod3a4 <= Co8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Vqd3a4 <= 1'b1;
	end
	else
	  begin
	    Vqd3a4 <= Mp8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Vsd3a4 <= 1'b0;
	end
	else
	  begin
	    Vsd3a4 <= Y78x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Wud3a4 <= 1'b1;
	end
	else
	  begin
	    Wud3a4 <= O07x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Swd3a4 <= 1'b1;
	end
	else
	  begin
	    Swd3a4 <= Joax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ryd3a4 <= 1'b0;
	end
	else
	  begin
	    Ryd3a4 <= Qb8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  S0e3a4 <= 1'b1;
	end
	else
	  begin
	    S0e3a4 <= Qw6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  P2e3a4 <= 1'b1;
	end
	else
	  begin
	    P2e3a4 <= Mmax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  P4e3a4 <= 1'b1;
	end
	else
	  begin
	    P4e3a4 <= Yy5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  P6e3a4 <= 1'b1;
	end
	else
	  begin
	    P6e3a4 <= My5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  P8e3a4 <= 1'b1;
	end
	else
	  begin
	    P8e3a4 <= Wk8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mae3a4 <= 1'b1;
	end
	else
	  begin
	    Mae3a4 <= Bkax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mce3a4 <= 1'b0;
	end
	else
	  begin
	    Mce3a4 <= Q88x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Lee3a4 <= 1'b0;
	end
	else
	  begin
	    Lee3a4 <= Gj8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Kge3a4 <= 1'b0;
	end
	else
	  begin
	    Kge3a4 <= Ad4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Iie3a4 <= 1'b1;
	end
	else
	  begin
	    Iie3a4 <= Sv7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hke3a4 <= 1'b0;
	end
	else
	  begin
	    Hke3a4 <= Uc4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Fme3a4 <= 1'b0;
	end
	else
	  begin
	    Fme3a4 <= Oc4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Doe3a4 <= 1'b0;
	end
	else
	  begin
	    Doe3a4 <= Lbax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Zpe3a4 <= 1'b0;
	end
	else
	  begin
	    Zpe3a4 <= Ncax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Vre3a4 <= 1'b1;
	end
	else
	  begin
	    Vre3a4 <= Sbax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rte3a4 <= 1'b0;
	end
	else
	  begin
	    Rte3a4 <= Uo8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Pve3a4 <= 1'b0;
	end
	else
	  begin
	    Pve3a4 <= Qw4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Jxe3a4 <= 1'b1;
	end
	else
	  begin
	    Jxe3a4 <= Kw4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Jze3a4 <= 1'b1;
	end
	else
	  begin
	    Jze3a4 <= Ic4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  G1f3a4 <= 1'b1;
	end
	else
	  begin
	    G1f3a4 <= Cc4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  G3f3a4 <= 1'b1;
	end
	else
	  begin
	    G3f3a4 <= Sm8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  G5f3a4 <= 1'b1;
	end
	else
	  begin
	    G5f3a4 <= Gs7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  F7f3a4 <= 1'b1;
	end
	else
	  begin
	    F7f3a4 <= O67x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  E9f3a4 <= 1'b1;
	end
	else
	  begin
	    E9f3a4 <= Q57x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Dbf3a4 <= 1'b1;
	end
	else
	  begin
	    Dbf3a4 <= Or6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Adf3a4 <= 1'b1;
	end
	else
	  begin
	    Adf3a4 <= U07x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xef3a4 <= 1'b1;
	end
	else
	  begin
	    Xef3a4 <= Gjax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xgf3a4 <= 1'b1;
	end
	else
	  begin
	    Xgf3a4 <= Ux4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xif3a4 <= 1'b1;
	end
	else
	  begin
	    Xif3a4 <= Ix4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xkf3a4 <= 1'b1;
	end
	else
	  begin
	    Xkf3a4 <= Kw6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Umf3a4 <= 1'b1;
	end
	else
	  begin
	    Umf3a4 <= Ikax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Uof3a4 <= 1'b1;
	end
	else
	  begin
	    Uof3a4 <= C95x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Uqf3a4 <= 1'b1;
	end
	else
	  begin
	    Uqf3a4 <= Q85x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Usf3a4 <= 1'b0;
	end
	else
	  begin
	    Usf3a4 <= Gcax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Quf3a4 <= 1'b0;
	end
	else
	  begin
	    Quf3a4 <= Wb4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rwf3a4 <= 1'b0;
	end
	else
	  begin
	    Rwf3a4 <= Ay7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Oyf3a4 <= 1'b1;
	end
	else
	  begin
	    Oyf3a4 <= K57x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  N0g3a4 <= 1'b1;
	end
	else
	  begin
	    N0g3a4 <= Ux6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  M2g3a4 <= 1'b1;
	end
	else
	  begin
	    M2g3a4 <= Ww6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  L4g3a4 <= 1'b1;
	end
	else
	  begin
	    L4g3a4 <= C08x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  I6g3a4 <= 1'b1;
	end
	else
	  begin
	    I6g3a4 <= Ujax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  I8g3a4 <= 1'b1;
	end
	else
	  begin
	    I8g3a4 <= E55x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Iag3a4 <= 1'b1;
	end
	else
	  begin
	    Iag3a4 <= S45x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Icg3a4 <= 1'b1;
	end
	else
	  begin
	    Icg3a4 <= Ma7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Heg3a4 <= 1'b0;
	end
	else
	  begin
	    Heg3a4 <= Oi8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hgg3a4 <= 1'b0;
	end
	else
	  begin
	    Hgg3a4 <= U98x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Jig3a4 <= 1'b1;
	end
	else
	  begin
	    Jig3a4 <= Ur8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ikg3a4 <= 1'b0;
	end
	else
	  begin
	    Ikg3a4 <= S48x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hmg3a4 <= 1'b0;
	end
	else
	  begin
	    Hmg3a4 <= Qb4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Gog3a4 <= 1'b0;
	end
	else
	  begin
	    Gog3a4 <= Aj8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Dqg3a4 <= 1'b0;
	end
	else
	  begin
	    Dqg3a4 <= Kb4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Csg3a4 <= 1'b1;
	end
	else
	  begin
	    Csg3a4 <= Eb4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cug3a4 <= 1'b1;
	end
	else
	  begin
	    Cug3a4 <= Ya4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cwg3a4 <= 1'b1;
	end
	else
	  begin
	    Cwg3a4 <= Sa4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cyg3a4 <= 1'b1;
	end
	else
	  begin
	    Cyg3a4 <= Ma4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  C0h3a4 <= 1'b1;
	end
	else
	  begin
	    C0h3a4 <= Ga4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  C2h3a4 <= 1'b1;
	end
	else
	  begin
	    C2h3a4 <= Aa4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  C4h3a4 <= 1'b1;
	end
	else
	  begin
	    C4h3a4 <= U94x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  B6h3a4 <= 1'b1;
	end
	else
	  begin
	    B6h3a4 <= O94x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  A8h3a4 <= 1'b1;
	end
	else
	  begin
	    A8h3a4 <= I94x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Z9h3a4 <= 1'b1;
	end
	else
	  begin
	    Z9h3a4 <= C94x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ybh3a4 <= 1'b1;
	end
	else
	  begin
	    Ybh3a4 <= W84x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xdh3a4 <= 1'b1;
	end
	else
	  begin
	    Xdh3a4 <= Q84x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Wfh3a4 <= 1'b1;
	end
	else
	  begin
	    Wfh3a4 <= K84x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Vhh3a4 <= 1'b1;
	end
	else
	  begin
	    Vhh3a4 <= E84x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ujh3a4 <= 1'b1;
	end
	else
	  begin
	    Ujh3a4 <= Y74x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Tlh3a4 <= 1'b1;
	end
	else
	  begin
	    Tlh3a4 <= S74x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Snh3a4 <= 1'b1;
	end
	else
	  begin
	    Snh3a4 <= Ap8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Sph3a4 <= 1'b1;
	end
	else
	  begin
	    Sph3a4 <= Ui8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Orh3a4 <= 1'b1;
	end
	else
	  begin
	    Orh3a4 <= M48x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Kth3a4 <= 1'b1;
	end
	else
	  begin
	    Kth3a4 <= O08x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Gvh3a4 <= 1'b1;
	end
	else
	  begin
	    Gvh3a4 <= Qz7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cxh3a4 <= 1'b1;
	end
	else
	  begin
	    Cxh3a4 <= Yy7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Yyh3a4 <= 1'b0;
	end
	else
	  begin
	    Yyh3a4 <= Nqax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  V0i3a4 <= 1'b1;
	end
	else
	  begin
	    V0i3a4 <= Ew6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  R2i3a4 <= 1'b1;
	end
	else
	  begin
	    R2i3a4 <= Ek4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  O4i3a4 <= 1'b1;
	end
	else
	  begin
	    O4i3a4 <= M74x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  L6i3a4 <= 1'b1;
	end
	else
	  begin
	    L6i3a4 <= G74x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  I8i3a4 <= 1'b1;
	end
	else
	  begin
	    I8i3a4 <= I38x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Iai3a4 <= 1'b1;
	end
	else
	  begin
	    Iai3a4 <= Y18x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hci3a4 <= 1'b1;
	end
	else
	  begin
	    Hci3a4 <= E28x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Gei3a4 <= 1'b1;
	end
	else
	  begin
	    Gei3a4 <= K28x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Fgi3a4 <= 1'b1;
	end
	else
	  begin
	    Fgi3a4 <= Q28x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Eii3a4 <= 1'b1;
	end
	else
	  begin
	    Eii3a4 <= W28x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Eki3a4 <= 1'b1;
	end
	else
	  begin
	    Eki3a4 <= C38x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Emi3a4 <= 1'b1;
	end
	else
	  begin
	    Emi3a4 <= O38x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Eoi3a4 <= 1'b1;
	end
	else
	  begin
	    Eoi3a4 <= U38x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Eqi3a4 <= 1'b1;
	end
	else
	  begin
	    Eqi3a4 <= Ym8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Esi3a4 <= 1'b1;
	end
	else
	  begin
	    Esi3a4 <= A48x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Eui3a4 <= 1'b1;
	end
	else
	  begin
	    Eui3a4 <= Zpax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Dwi3a4 <= 1'b1;
	end
	else
	  begin
	    Dwi3a4 <= S18x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cyi3a4 <= 1'b0;
	end
	else
	  begin
	    Cyi3a4 <= Ux7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Zzi3a4 <= 1'b1;
	end
	else
	  begin
	    Zzi3a4 <= Mv7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Y1j3a4 <= 1'b1;
	end
	else
	  begin
	    Y1j3a4 <= Yv7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  X3j3a4 <= 1'b1;
	end
	else
	  begin
	    X3j3a4 <= Ew7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  W5j3a4 <= 1'b1;
	end
	else
	  begin
	    W5j3a4 <= Kw7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  V7j3a4 <= 1'b1;
	end
	else
	  begin
	    V7j3a4 <= Qw7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  U9j3a4 <= 1'b1;
	end
	else
	  begin
	    U9j3a4 <= Ww7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ubj3a4 <= 1'b1;
	end
	else
	  begin
	    Ubj3a4 <= Cx7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Udj3a4 <= 1'b1;
	end
	else
	  begin
	    Udj3a4 <= Ix7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ufj3a4 <= 1'b0;
	end
	else
	  begin
	    Ufj3a4 <= Gv7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rhj3a4 <= 1'b1;
	end
	else
	  begin
	    Rhj3a4 <= Ox7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rjj3a4 <= 1'b1;
	end
	else
	  begin
	    Rjj3a4 <= K58x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Qlj3a4 <= 1'b1;
	end
	else
	  begin
	    Qlj3a4 <= Oo8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Qnj3a4 <= 1'b1;
	end
	else
	  begin
	    Qnj3a4 <= Ss8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Tpj3a4 <= 1'b1;
	end
	else
	  begin
	    Tpj3a4 <= Ir8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Srj3a4 <= 1'b1;
	end
	else
	  begin
	    Srj3a4 <= Or8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rtj3a4 <= 1'b1;
	end
	else
	  begin
	    Rtj3a4 <= Kt7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Qvj3a4 <= 1'b1;
	end
	else
	  begin
	    Qvj3a4 <= Qt7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Pxj3a4 <= 1'b1;
	end
	else
	  begin
	    Pxj3a4 <= Wt7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ozj3a4 <= 1'b1;
	end
	else
	  begin
	    Ozj3a4 <= Yp8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  N1k3a4 <= 1'b1;
	end
	else
	  begin
	    N1k3a4 <= Ur7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  M3k3a4 <= 1'b1;
	end
	else
	  begin
	    M3k3a4 <= Ii7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  M5k3a4 <= 1'b1;
	end
	else
	  begin
	    M5k3a4 <= Qh7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  L7k3a4 <= 1'b1;
	end
	else
	  begin
	    L7k3a4 <= W87x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  K9k3a4 <= 1'b1;
	end
	else
	  begin
	    K9k3a4 <= Y47x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Jbk3a4 <= 1'b1;
	end
	else
	  begin
	    Jbk3a4 <= C07x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Idk3a4 <= 1'b1;
	end
	else
	  begin
	    Idk3a4 <= Mv6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hfk3a4 <= 1'b1;
	end
	else
	  begin
	    Hfk3a4 <= Cr6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ghk3a4 <= 1'b1;
	end
	else
	  begin
	    Ghk3a4 <= Ag6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Fjk3a4 <= 1'b1;
	end
	else
	  begin
	    Fjk3a4 <= G16x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Flk3a4 <= 1'b1;
	end
	else
	  begin
	    Flk3a4 <= Ox5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Fnk3a4 <= 1'b1;
	end
	else
	  begin
	    Fnk3a4 <= Wt5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Fpk3a4 <= 1'b1;
	end
	else
	  begin
	    Fpk3a4 <= Ui5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Frk3a4 <= 1'b1;
	end
	else
	  begin
	    Frk3a4 <= Kb5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ftk3a4 <= 1'b1;
	end
	else
	  begin
	    Ftk3a4 <= M75x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Fvk3a4 <= 1'b1;
	end
	else
	  begin
	    Fvk3a4 <= U35x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Fxk3a4 <= 1'b1;
	end
	else
	  begin
	    Fxk3a4 <= C05x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Fzk3a4 <= 1'b1;
	end
	else
	  begin
	    Fzk3a4 <= Yv4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  F1l3a4 <= 1'b1;
	end
	else
	  begin
	    F1l3a4 <= Ur4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  F3l3a4 <= 1'b1;
	end
	else
	  begin
	    F3l3a4 <= Qn4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  F5l3a4 <= 1'b1;
	end
	else
	  begin
	    F5l3a4 <= Mj4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  F7l3a4 <= 1'b1;
	end
	else
	  begin
	    F7l3a4 <= Qk7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  E9l3a4 <= 1'b1;
	end
	else
	  begin
	    E9l3a4 <= Kk7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Dbl3a4 <= 1'b1;
	end
	else
	  begin
	    Dbl3a4 <= Ek7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cdl3a4 <= 1'b1;
	end
	else
	  begin
	    Cdl3a4 <= Mj7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cfl3a4 <= 1'b1;
	end
	else
	  begin
	    Cfl3a4 <= E87x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Bhl3a4 <= 1'b1;
	end
	else
	  begin
	    Bhl3a4 <= G47x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ajl3a4 <= 1'b1;
	end
	else
	  begin
	    Ajl3a4 <= Kz6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Zkl3a4 <= 1'b1;
	end
	else
	  begin
	    Zkl3a4 <= Uu6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Yml3a4 <= 1'b1;
	end
	else
	  begin
	    Yml3a4 <= Kq6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xol3a4 <= 1'b1;
	end
	else
	  begin
	    Xol3a4 <= If6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xql3a4 <= 1'b1;
	end
	else
	  begin
	    Xql3a4 <= O06x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xsl3a4 <= 1'b1;
	end
	else
	  begin
	    Xsl3a4 <= Ww5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xul3a4 <= 1'b1;
	end
	else
	  begin
	    Xul3a4 <= Et5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xwl3a4 <= 1'b1;
	end
	else
	  begin
	    Xwl3a4 <= Ci5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xyl3a4 <= 1'b1;
	end
	else
	  begin
	    Xyl3a4 <= Sa5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  X0m3a4 <= 1'b1;
	end
	else
	  begin
	    X0m3a4 <= U65x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  X2m3a4 <= 1'b1;
	end
	else
	  begin
	    X2m3a4 <= C35x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  X4m3a4 <= 1'b1;
	end
	else
	  begin
	    X4m3a4 <= Kz4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  X6m3a4 <= 1'b1;
	end
	else
	  begin
	    X6m3a4 <= Gv4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  X8m3a4 <= 1'b1;
	end
	else
	  begin
	    X8m3a4 <= Cr4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xam3a4 <= 1'b1;
	end
	else
	  begin
	    Xam3a4 <= Ym4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xcm3a4 <= 1'b1;
	end
	else
	  begin
	    Xcm3a4 <= Ui4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xem3a4 <= 1'b1;
	end
	else
	  begin
	    Xem3a4 <= Oi4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xgm3a4 <= 1'b1;
	end
	else
	  begin
	    Xgm3a4 <= Sm4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xim3a4 <= 1'b1;
	end
	else
	  begin
	    Xim3a4 <= Wq4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xkm3a4 <= 1'b1;
	end
	else
	  begin
	    Xkm3a4 <= Av4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xmm3a4 <= 1'b1;
	end
	else
	  begin
	    Xmm3a4 <= Ez4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xom3a4 <= 1'b1;
	end
	else
	  begin
	    Xom3a4 <= W25x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xqm3a4 <= 1'b1;
	end
	else
	  begin
	    Xqm3a4 <= O65x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xsm3a4 <= 1'b1;
	end
	else
	  begin
	    Xsm3a4 <= Ma5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xum3a4 <= 1'b1;
	end
	else
	  begin
	    Xum3a4 <= Wh5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xwm3a4 <= 1'b1;
	end
	else
	  begin
	    Xwm3a4 <= Ys5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xym3a4 <= 1'b1;
	end
	else
	  begin
	    Xym3a4 <= Qw5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  X0n3a4 <= 1'b1;
	end
	else
	  begin
	    X0n3a4 <= I06x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  X2n3a4 <= 1'b1;
	end
	else
	  begin
	    X2n3a4 <= Cf6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  X4n3a4 <= 1'b1;
	end
	else
	  begin
	    X4n3a4 <= Eq6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  W6n3a4 <= 1'b1;
	end
	else
	  begin
	    W6n3a4 <= Ou6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  V8n3a4 <= 1'b1;
	end
	else
	  begin
	    V8n3a4 <= Ez6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Uan3a4 <= 1'b1;
	end
	else
	  begin
	    Uan3a4 <= A47x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Tcn3a4 <= 1'b1;
	end
	else
	  begin
	    Tcn3a4 <= Y77x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Sen3a4 <= 1'b1;
	end
	else
	  begin
	    Sen3a4 <= Wk7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Sgn3a4 <= 1'b1;
	end
	else
	  begin
	    Sgn3a4 <= Ol7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rin3a4 <= 1'b1;
	end
	else
	  begin
	    Rin3a4 <= Ul7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Qkn3a4 <= 1'b1;
	end
	else
	  begin
	    Qkn3a4 <= Am7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Pmn3a4 <= 1'b1;
	end
	else
	  begin
	    Pmn3a4 <= Kn7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Oon3a4 <= 1'b1;
	end
	else
	  begin
	    Oon3a4 <= En7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Nqn3a4 <= 1'b1;
	end
	else
	  begin
	    Nqn3a4 <= Ym7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Msn3a4 <= 1'b1;
	end
	else
	  begin
	    Msn3a4 <= Gm7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mun3a4 <= 1'b1;
	end
	else
	  begin
	    Mun3a4 <= S77x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Lwn3a4 <= 1'b1;
	end
	else
	  begin
	    Lwn3a4 <= U37x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Kyn3a4 <= 1'b1;
	end
	else
	  begin
	    Kyn3a4 <= Yy6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  J0o3a4 <= 1'b1;
	end
	else
	  begin
	    J0o3a4 <= Iu6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  I2o3a4 <= 1'b1;
	end
	else
	  begin
	    I2o3a4 <= Yp6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  H4o3a4 <= 1'b1;
	end
	else
	  begin
	    H4o3a4 <= We6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  H6o3a4 <= 1'b1;
	end
	else
	  begin
	    H6o3a4 <= C06x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  H8o3a4 <= 1'b1;
	end
	else
	  begin
	    H8o3a4 <= Kw5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hao3a4 <= 1'b1;
	end
	else
	  begin
	    Hao3a4 <= Ss5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hco3a4 <= 1'b1;
	end
	else
	  begin
	    Hco3a4 <= Qh5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Heo3a4 <= 1'b1;
	end
	else
	  begin
	    Heo3a4 <= Ga5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hgo3a4 <= 1'b1;
	end
	else
	  begin
	    Hgo3a4 <= I65x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hio3a4 <= 1'b1;
	end
	else
	  begin
	    Hio3a4 <= Q25x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hko3a4 <= 1'b1;
	end
	else
	  begin
	    Hko3a4 <= Yy4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hmo3a4 <= 1'b1;
	end
	else
	  begin
	    Hmo3a4 <= Uu4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hoo3a4 <= 1'b1;
	end
	else
	  begin
	    Hoo3a4 <= Qq4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hqo3a4 <= 1'b1;
	end
	else
	  begin
	    Hqo3a4 <= Mm4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hso3a4 <= 1'b1;
	end
	else
	  begin
	    Hso3a4 <= Ii4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Huo3a4 <= 1'b1;
	end
	else
	  begin
	    Huo3a4 <= Ci4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hwo3a4 <= 1'b1;
	end
	else
	  begin
	    Hwo3a4 <= Gm4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hyo3a4 <= 1'b1;
	end
	else
	  begin
	    Hyo3a4 <= Kq4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  H0p3a4 <= 1'b1;
	end
	else
	  begin
	    H0p3a4 <= Ou4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  H2p3a4 <= 1'b1;
	end
	else
	  begin
	    H2p3a4 <= Sy4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  H4p3a4 <= 1'b1;
	end
	else
	  begin
	    H4p3a4 <= K25x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  H6p3a4 <= 1'b1;
	end
	else
	  begin
	    H6p3a4 <= C65x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  H8p3a4 <= 1'b1;
	end
	else
	  begin
	    H8p3a4 <= Aa5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hap3a4 <= 1'b1;
	end
	else
	  begin
	    Hap3a4 <= Kh5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hcp3a4 <= 1'b1;
	end
	else
	  begin
	    Hcp3a4 <= Ms5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hep3a4 <= 1'b1;
	end
	else
	  begin
	    Hep3a4 <= Ew5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hgp3a4 <= 1'b1;
	end
	else
	  begin
	    Hgp3a4 <= Wz5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hip3a4 <= 1'b1;
	end
	else
	  begin
	    Hip3a4 <= Qe6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hkp3a4 <= 1'b1;
	end
	else
	  begin
	    Hkp3a4 <= Sp6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Gmp3a4 <= 1'b1;
	end
	else
	  begin
	    Gmp3a4 <= Cu6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Fop3a4 <= 1'b1;
	end
	else
	  begin
	    Fop3a4 <= Sy6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Eqp3a4 <= 1'b1;
	end
	else
	  begin
	    Eqp3a4 <= O37x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Dsp3a4 <= 1'b1;
	end
	else
	  begin
	    Dsp3a4 <= M77x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cup3a4 <= 1'b1;
	end
	else
	  begin
	    Cup3a4 <= Qn7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cwp3a4 <= 1'b1;
	end
	else
	  begin
	    Cwp3a4 <= Io7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Byp3a4 <= 1'b1;
	end
	else
	  begin
	    Byp3a4 <= Oo7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  A0q3a4 <= 1'b1;
	end
	else
	  begin
	    A0q3a4 <= Uo7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Z1q3a4 <= 1'b1;
	end
	else
	  begin
	    Z1q3a4 <= Eq7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Y3q3a4 <= 1'b1;
	end
	else
	  begin
	    Y3q3a4 <= Yp7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  X5q3a4 <= 1'b1;
	end
	else
	  begin
	    X5q3a4 <= Sp7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  W7q3a4 <= 1'b1;
	end
	else
	  begin
	    W7q3a4 <= Ap7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  W9q3a4 <= 1'b1;
	end
	else
	  begin
	    W9q3a4 <= I67x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Vbq3a4 <= 1'b1;
	end
	else
	  begin
	    Vbq3a4 <= K27x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Udq3a4 <= 1'b1;
	end
	else
	  begin
	    Udq3a4 <= Ox6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Tfq3a4 <= 1'b1;
	end
	else
	  begin
	    Tfq3a4 <= Ys6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Shq3a4 <= 1'b1;
	end
	else
	  begin
	    Shq3a4 <= Oo6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rjq3a4 <= 1'b1;
	end
	else
	  begin
	    Rjq3a4 <= Md6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rlq3a4 <= 1'b1;
	end
	else
	  begin
	    Rlq3a4 <= Sy5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rnq3a4 <= 1'b1;
	end
	else
	  begin
	    Rnq3a4 <= Av5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rpq3a4 <= 1'b1;
	end
	else
	  begin
	    Rpq3a4 <= Ir5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rrq3a4 <= 1'b1;
	end
	else
	  begin
	    Rrq3a4 <= Gg5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rtq3a4 <= 1'b1;
	end
	else
	  begin
	    Rtq3a4 <= W85x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rvq3a4 <= 1'b1;
	end
	else
	  begin
	    Rvq3a4 <= Y45x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rxq3a4 <= 1'b1;
	end
	else
	  begin
	    Rxq3a4 <= G15x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rzq3a4 <= 1'b1;
	end
	else
	  begin
	    Rzq3a4 <= Ox4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  R1r3a4 <= 1'b1;
	end
	else
	  begin
	    R1r3a4 <= Kt4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  R3r3a4 <= 1'b1;
	end
	else
	  begin
	    R3r3a4 <= Gp4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  R5r3a4 <= 1'b1;
	end
	else
	  begin
	    R5r3a4 <= Cl4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  R7r3a4 <= 1'b1;
	end
	else
	  begin
	    R7r3a4 <= Yg4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  R9r3a4 <= 1'b1;
	end
	else
	  begin
	    R9r3a4 <= Or7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Qbr3a4 <= 1'b1;
	end
	else
	  begin
	    Qbr3a4 <= Ir7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Pdr3a4 <= 1'b1;
	end
	else
	  begin
	    Pdr3a4 <= Cr7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ofr3a4 <= 1'b1;
	end
	else
	  begin
	    Ofr3a4 <= Kq7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ohr3a4 <= 1'b1;
	end
	else
	  begin
	    Ohr3a4 <= W57x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Njr3a4 <= 1'b1;
	end
	else
	  begin
	    Njr3a4 <= Y17x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mlr3a4 <= 1'b1;
	end
	else
	  begin
	    Mlr3a4 <= Cx6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Lnr3a4 <= 1'b1;
	end
	else
	  begin
	    Lnr3a4 <= Ms6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Kpr3a4 <= 1'b1;
	end
	else
	  begin
	    Kpr3a4 <= Io6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Jrr3a4 <= 1'b1;
	end
	else
	  begin
	    Jrr3a4 <= Cr5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Jtr3a4 <= 1'b1;
	end
	else
	  begin
	    Jtr3a4 <= Et4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Jvr3a4 <= 1'b1;
	end
	else
	  begin
	    Jvr3a4 <= Ap4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Jxr3a4 <= 1'b1;
	end
	else
	  begin
	    Jxr3a4 <= Mg4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Jzr3a4 <= 1'b1;
	end
	else
	  begin
	    Jzr3a4 <= Sg4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  J1s3a4 <= 1'b1;
	end
	else
	  begin
	    J1s3a4 <= Wk4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  J3s3a4 <= 1'b1;
	end
	else
	  begin
	    J3s3a4 <= Ss4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  J5s3a4 <= 1'b1;
	end
	else
	  begin
	    J5s3a4 <= Ww4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  J7s3a4 <= 1'b1;
	end
	else
	  begin
	    J7s3a4 <= O05x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  J9s3a4 <= 1'b1;
	end
	else
	  begin
	    J9s3a4 <= G45x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Jbs3a4 <= 1'b1;
	end
	else
	  begin
	    Jbs3a4 <= Y75x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Jds3a4 <= 1'b1;
	end
	else
	  begin
	    Jds3a4 <= Wb5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Jfs3a4 <= 1'b1;
	end
	else
	  begin
	    Jfs3a4 <= Gj5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Jhs3a4 <= 1'b1;
	end
	else
	  begin
	    Jhs3a4 <= Ay5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Jjs3a4 <= 1'b1;
	end
	else
	  begin
	    Jjs3a4 <= S16x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Jls3a4 <= 1'b1;
	end
	else
	  begin
	    Jls3a4 <= Mg6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Jns3a4 <= 1'b1;
	end
	else
	  begin
	    Jns3a4 <= Ss6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ips3a4 <= 1'b1;
	end
	else
	  begin
	    Ips3a4 <= Ix6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hrs3a4 <= 1'b1;
	end
	else
	  begin
	    Hrs3a4 <= E27x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Gts3a4 <= 1'b1;
	end
	else
	  begin
	    Gts3a4 <= C67x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Fvs3a4 <= 1'b1;
	end
	else
	  begin
	    Fvs3a4 <= I68x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Exs3a4 <= 1'b1;
	end
	else
	  begin
	    Exs3a4 <= O68x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Dzs3a4 <= 1'b1;
	end
	else
	  begin
	    Dzs3a4 <= U68x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  C1t3a4 <= 1'b1;
	end
	else
	  begin
	    C1t3a4 <= Iu5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  C3t3a4 <= 1'b1;
	end
	else
	  begin
	    C3t3a4 <= Gg4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  C5t3a4 <= 1'b1;
	end
	else
	  begin
	    C5t3a4 <= Kk4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  C7t3a4 <= 1'b1;
	end
	else
	  begin
	    C7t3a4 <= Cx4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  C9t3a4 <= 1'b1;
	end
	else
	  begin
	    C9t3a4 <= U05x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cbt3a4 <= 1'b1;
	end
	else
	  begin
	    Cbt3a4 <= M45x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cdt3a4 <= 1'b1;
	end
	else
	  begin
	    Cdt3a4 <= K85x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cft3a4 <= 1'b1;
	end
	else
	  begin
	    Cft3a4 <= Uf5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cht3a4 <= 1'b1;
	end
	else
	  begin
	    Cht3a4 <= Ou5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cjt3a4 <= 1'b1;
	end
	else
	  begin
	    Cjt3a4 <= Gy5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Clt3a4 <= 1'b1;
	end
	else
	  begin
	    Clt3a4 <= Ad6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cnt3a4 <= 1'b1;
	end
	else
	  begin
	    Cnt3a4 <= Co6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Bpt3a4 <= 1'b1;
	end
	else
	  begin
	    Bpt3a4 <= M78x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Art3a4 <= 1'b1;
	end
	else
	  begin
	    Art3a4 <= Ol8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Zst3a4 <= 1'b1;
	end
	else
	  begin
	    Zst3a4 <= Ul8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Zut3a4 <= 1'b1;
	end
	else
	  begin
	    Zut3a4 <= Gj7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Zwt3a4 <= 1'b1;
	end
	else
	  begin
	    Zwt3a4 <= Oi7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Yyt3a4 <= 1'b1;
	end
	else
	  begin
	    Yyt3a4 <= C97x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  X0u3a4 <= 1'b1;
	end
	else
	  begin
	    X0u3a4 <= E57x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  W2u3a4 <= 1'b1;
	end
	else
	  begin
	    W2u3a4 <= I07x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  V4u3a4 <= 1'b1;
	end
	else
	  begin
	    V4u3a4 <= Sv6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  U6u3a4 <= 1'b1;
	end
	else
	  begin
	    U6u3a4 <= Ir6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  T8u3a4 <= 1'b1;
	end
	else
	  begin
	    T8u3a4 <= Gg6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Sau3a4 <= 1'b1;
	end
	else
	  begin
	    Sau3a4 <= M16x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Scu3a4 <= 1'b1;
	end
	else
	  begin
	    Scu3a4 <= Ux5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Seu3a4 <= 1'b1;
	end
	else
	  begin
	    Seu3a4 <= Cu5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Sgu3a4 <= 1'b1;
	end
	else
	  begin
	    Sgu3a4 <= Aj5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Siu3a4 <= 1'b1;
	end
	else
	  begin
	    Siu3a4 <= Qb5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Sku3a4 <= 1'b1;
	end
	else
	  begin
	    Sku3a4 <= S75x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Smu3a4 <= 1'b1;
	end
	else
	  begin
	    Smu3a4 <= A45x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Sou3a4 <= 1'b1;
	end
	else
	  begin
	    Sou3a4 <= I05x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Squ3a4 <= 1'b1;
	end
	else
	  begin
	    Squ3a4 <= Ew4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ssu3a4 <= 1'b1;
	end
	else
	  begin
	    Ssu3a4 <= As4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Suu3a4 <= 1'b1;
	end
	else
	  begin
	    Suu3a4 <= Wn4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Swu3a4 <= 1'b1;
	end
	else
	  begin
	    Swu3a4 <= Sj4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Syu3a4 <= 1'b1;
	end
	else
	  begin
	    Syu3a4 <= Kh7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  R0v3a4 <= 1'b1;
	end
	else
	  begin
	    R0v3a4 <= Eh7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Q2v3a4 <= 1'b1;
	end
	else
	  begin
	    Q2v3a4 <= Yg7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  P4v3a4 <= 1'b1;
	end
	else
	  begin
	    P4v3a4 <= Gg7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  P6v3a4 <= 1'b1;
	end
	else
	  begin
	    P6v3a4 <= Q87x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  O8v3a4 <= 1'b1;
	end
	else
	  begin
	    O8v3a4 <= S47x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Nav3a4 <= 1'b1;
	end
	else
	  begin
	    Nav3a4 <= Wz6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mcv3a4 <= 1'b1;
	end
	else
	  begin
	    Mcv3a4 <= Gv6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Lev3a4 <= 1'b1;
	end
	else
	  begin
	    Lev3a4 <= Wq6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Kgv3a4 <= 1'b1;
	end
	else
	  begin
	    Kgv3a4 <= Uf6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Kiv3a4 <= 1'b1;
	end
	else
	  begin
	    Kiv3a4 <= A16x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Kkv3a4 <= 1'b1;
	end
	else
	  begin
	    Kkv3a4 <= Ix5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Kmv3a4 <= 1'b1;
	end
	else
	  begin
	    Kmv3a4 <= Qt5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Kov3a4 <= 1'b1;
	end
	else
	  begin
	    Kov3a4 <= Oi5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Kqv3a4 <= 1'b1;
	end
	else
	  begin
	    Kqv3a4 <= Eb5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ksv3a4 <= 1'b1;
	end
	else
	  begin
	    Ksv3a4 <= G75x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Kuv3a4 <= 1'b1;
	end
	else
	  begin
	    Kuv3a4 <= O35x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Kwv3a4 <= 1'b1;
	end
	else
	  begin
	    Kwv3a4 <= Wz4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Kyv3a4 <= 1'b1;
	end
	else
	  begin
	    Kyv3a4 <= Sv4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  K0w3a4 <= 1'b1;
	end
	else
	  begin
	    K0w3a4 <= Or4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  K2w3a4 <= 1'b1;
	end
	else
	  begin
	    K2w3a4 <= Kn4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  K4w3a4 <= 1'b1;
	end
	else
	  begin
	    K4w3a4 <= Gj4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  K6w3a4 <= 1'b1;
	end
	else
	  begin
	    K6w3a4 <= Ag7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  J8w3a4 <= 1'b1;
	end
	else
	  begin
	    J8w3a4 <= Uf7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Iaw3a4 <= 1'b1;
	end
	else
	  begin
	    Iaw3a4 <= Of7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hcw3a4 <= 1'b1;
	end
	else
	  begin
	    Hcw3a4 <= We7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hew3a4 <= 1'b1;
	end
	else
	  begin
	    Hew3a4 <= K87x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ggw3a4 <= 1'b1;
	end
	else
	  begin
	    Ggw3a4 <= M47x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Fiw3a4 <= 1'b1;
	end
	else
	  begin
	    Fiw3a4 <= Qz6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ekw3a4 <= 1'b1;
	end
	else
	  begin
	    Ekw3a4 <= Av6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Dmw3a4 <= 1'b1;
	end
	else
	  begin
	    Dmw3a4 <= Qq6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cow3a4 <= 1'b1;
	end
	else
	  begin
	    Cow3a4 <= Of6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cqw3a4 <= 1'b1;
	end
	else
	  begin
	    Cqw3a4 <= U06x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Csw3a4 <= 1'b1;
	end
	else
	  begin
	    Csw3a4 <= Cx5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cuw3a4 <= 1'b1;
	end
	else
	  begin
	    Cuw3a4 <= Kt5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cww3a4 <= 1'b1;
	end
	else
	  begin
	    Cww3a4 <= Ii5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cyw3a4 <= 1'b1;
	end
	else
	  begin
	    Cyw3a4 <= Ya5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  C0x3a4 <= 1'b1;
	end
	else
	  begin
	    C0x3a4 <= A75x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  C2x3a4 <= 1'b1;
	end
	else
	  begin
	    C2x3a4 <= I35x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  C4x3a4 <= 1'b1;
	end
	else
	  begin
	    C4x3a4 <= Qz4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  C6x3a4 <= 1'b1;
	end
	else
	  begin
	    C6x3a4 <= Mv4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  C8x3a4 <= 1'b1;
	end
	else
	  begin
	    C8x3a4 <= Ir4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cax3a4 <= 1'b1;
	end
	else
	  begin
	    Cax3a4 <= En4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ccx3a4 <= 1'b1;
	end
	else
	  begin
	    Ccx3a4 <= Aj4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cex3a4 <= 1'b1;
	end
	else
	  begin
	    Cex3a4 <= Wb7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Bgx3a4 <= 1'b1;
	end
	else
	  begin
	    Bgx3a4 <= Qb7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Aix3a4 <= 1'b1;
	end
	else
	  begin
	    Aix3a4 <= Kb7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Zjx3a4 <= 1'b1;
	end
	else
	  begin
	    Zjx3a4 <= Sa7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Zlx3a4 <= 1'b1;
	end
	else
	  begin
	    Zlx3a4 <= U67x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ynx3a4 <= 1'b1;
	end
	else
	  begin
	    Ynx3a4 <= W27x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xpx3a4 <= 1'b1;
	end
	else
	  begin
	    Xpx3a4 <= Ay6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Wrx3a4 <= 1'b1;
	end
	else
	  begin
	    Wrx3a4 <= Kt6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Vtx3a4 <= 1'b1;
	end
	else
	  begin
	    Vtx3a4 <= Ap6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Uvx3a4 <= 1'b1;
	end
	else
	  begin
	    Uvx3a4 <= Yd6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Uxx3a4 <= 1'b1;
	end
	else
	  begin
	    Uxx3a4 <= Ez5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Uzx3a4 <= 1'b1;
	end
	else
	  begin
	    Uzx3a4 <= Mv5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  U1y3a4 <= 1'b1;
	end
	else
	  begin
	    U1y3a4 <= Ur5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  U3y3a4 <= 1'b1;
	end
	else
	  begin
	    U3y3a4 <= Sg5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  U5y3a4 <= 1'b1;
	end
	else
	  begin
	    U5y3a4 <= I95x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  U7y3a4 <= 1'b1;
	end
	else
	  begin
	    U7y3a4 <= K55x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  U9y3a4 <= 1'b1;
	end
	else
	  begin
	    U9y3a4 <= S15x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Uby3a4 <= 1'b1;
	end
	else
	  begin
	    Uby3a4 <= Ay4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Udy3a4 <= 1'b1;
	end
	else
	  begin
	    Udy3a4 <= Wt4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ufy3a4 <= 1'b1;
	end
	else
	  begin
	    Ufy3a4 <= Sp4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Uhy3a4 <= 1'b1;
	end
	else
	  begin
	    Uhy3a4 <= Ol4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ujy3a4 <= 1'b1;
	end
	else
	  begin
	    Ujy3a4 <= Kh4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Uly3a4 <= 1'b1;
	end
	else
	  begin
	    Uly3a4 <= Gd7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Tny3a4 <= 1'b1;
	end
	else
	  begin
	    Tny3a4 <= Ad7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Spy3a4 <= 1'b1;
	end
	else
	  begin
	    Spy3a4 <= Uc7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rry3a4 <= 1'b1;
	end
	else
	  begin
	    Rry3a4 <= Cc7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rty3a4 <= 1'b1;
	end
	else
	  begin
	    Rty3a4 <= A77x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Qvy3a4 <= 1'b1;
	end
	else
	  begin
	    Qvy3a4 <= C37x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Pxy3a4 <= 1'b1;
	end
	else
	  begin
	    Pxy3a4 <= Gy6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ozy3a4 <= 1'b1;
	end
	else
	  begin
	    Ozy3a4 <= Qt6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  N1z3a4 <= 1'b1;
	end
	else
	  begin
	    N1z3a4 <= Gp6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  M3z3a4 <= 1'b1;
	end
	else
	  begin
	    M3z3a4 <= Ee6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  M5z3a4 <= 1'b1;
	end
	else
	  begin
	    M5z3a4 <= Kz5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  M7z3a4 <= 1'b1;
	end
	else
	  begin
	    M7z3a4 <= Sv5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  M9z3a4 <= 1'b1;
	end
	else
	  begin
	    M9z3a4 <= As5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mbz3a4 <= 1'b1;
	end
	else
	  begin
	    Mbz3a4 <= Yg5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mdz3a4 <= 1'b1;
	end
	else
	  begin
	    Mdz3a4 <= O95x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mfz3a4 <= 1'b1;
	end
	else
	  begin
	    Mfz3a4 <= Q55x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mhz3a4 <= 1'b1;
	end
	else
	  begin
	    Mhz3a4 <= Y15x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mjz3a4 <= 1'b1;
	end
	else
	  begin
	    Mjz3a4 <= Gy4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mlz3a4 <= 1'b1;
	end
	else
	  begin
	    Mlz3a4 <= Cu4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mnz3a4 <= 1'b1;
	end
	else
	  begin
	    Mnz3a4 <= Yp4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mpz3a4 <= 1'b1;
	end
	else
	  begin
	    Mpz3a4 <= Ul4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mrz3a4 <= 1'b1;
	end
	else
	  begin
	    Mrz3a4 <= Qh4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mtz3a4 <= 1'b1;
	end
	else
	  begin
	    Mtz3a4 <= Wh4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mvz3a4 <= 1'b1;
	end
	else
	  begin
	    Mvz3a4 <= Am4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mxz3a4 <= 1'b1;
	end
	else
	  begin
	    Mxz3a4 <= Eq4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mzz3a4 <= 1'b1;
	end
	else
	  begin
	    Mzz3a4 <= Iu4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  M104a4 <= 1'b1;
	end
	else
	  begin
	    M104a4 <= My4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  M304a4 <= 1'b1;
	end
	else
	  begin
	    M304a4 <= E25x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  M504a4 <= 1'b1;
	end
	else
	  begin
	    M504a4 <= W55x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  M704a4 <= 1'b1;
	end
	else
	  begin
	    M704a4 <= U95x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  M904a4 <= 1'b1;
	end
	else
	  begin
	    M904a4 <= Eh5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mb04a4 <= 1'b1;
	end
	else
	  begin
	    Mb04a4 <= Gs5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Md04a4 <= 1'b1;
	end
	else
	  begin
	    Md04a4 <= Yv5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mf04a4 <= 1'b1;
	end
	else
	  begin
	    Mf04a4 <= Qz5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mh04a4 <= 1'b1;
	end
	else
	  begin
	    Mh04a4 <= Sa6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mj04a4 <= 1'b1;
	end
	else
	  begin
	    Mj04a4 <= I96x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ml04a4 <= 1'b1;
	end
	else
	  begin
	    Ml04a4 <= Ya6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mn04a4 <= 1'b1;
	end
	else
	  begin
	    Mn04a4 <= Kb6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mp04a4 <= 1'b1;
	end
	else
	  begin
	    Mp04a4 <= Uc6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mr04a4 <= 1'b1;
	end
	else
	  begin
	    Mr04a4 <= Oc6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Lt04a4 <= 1'b1;
	end
	else
	  begin
	    Lt04a4 <= Ic6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Kv04a4 <= 1'b1;
	end
	else
	  begin
	    Kv04a4 <= Cc6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Kx04a4 <= 1'b1;
	end
	else
	  begin
	    Kx04a4 <= Wb6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Kz04a4 <= 1'b1;
	end
	else
	  begin
	    Kz04a4 <= Qb6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  K114a4 <= 1'b1;
	end
	else
	  begin
	    K114a4 <= Eb6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  K314a4 <= 1'b1;
	end
	else
	  begin
	    K314a4 <= Ma6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  K514a4 <= 1'b1;
	end
	else
	  begin
	    K514a4 <= Ga6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  K714a4 <= 1'b1;
	end
	else
	  begin
	    K714a4 <= Aa6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  K914a4 <= 1'b1;
	end
	else
	  begin
	    K914a4 <= U96x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Kb14a4 <= 1'b1;
	end
	else
	  begin
	    Kb14a4 <= O96x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Kd14a4 <= 1'b1;
	end
	else
	  begin
	    Kd14a4 <= Ke6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Kf14a4 <= 1'b1;
	end
	else
	  begin
	    Kf14a4 <= Wt6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Jh14a4 <= 1'b1;
	end
	else
	  begin
	    Jh14a4 <= My6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ij14a4 <= 1'b1;
	end
	else
	  begin
	    Ij14a4 <= I37x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hl14a4 <= 1'b1;
	end
	else
	  begin
	    Hl14a4 <= G77x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Gn14a4 <= 1'b1;
	end
	else
	  begin
	    Gn14a4 <= Md7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Gp14a4 <= 1'b1;
	end
	else
	  begin
	    Gp14a4 <= Yd7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Gr14a4 <= 1'b1;
	end
	else
	  begin
	    Gr14a4 <= E85x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Gt14a4 <= 1'b1;
	end
	else
	  begin
	    Gt14a4 <= Wh7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Gv14a4 <= 1'b1;
	end
	else
	  begin
	    Gv14a4 <= Il7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Gx14a4 <= 1'b1;
	end
	else
	  begin
	    Gx14a4 <= Co7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Gz14a4 <= 1'b1;
	end
	else
	  begin
	    Gz14a4 <= Qk8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  G124a4 <= 1'b1;
	end
	else
	  begin
	    G124a4 <= Wq7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  G324a4 <= 1'b1;
	end
	else
	  begin
	    G324a4 <= Mp7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  G524a4 <= 1'b1;
	end
	else
	  begin
	    G524a4 <= Sm7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  G724a4 <= 1'b1;
	end
	else
	  begin
	    G724a4 <= Yj7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  G924a4 <= 1'b1;
	end
	else
	  begin
	    G924a4 <= Ui7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Gb24a4 <= 1'b1;
	end
	else
	  begin
	    Gb24a4 <= Sg7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Gd24a4 <= 1'b1;
	end
	else
	  begin
	    Gd24a4 <= If7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Gf24a4 <= 1'b1;
	end
	else
	  begin
	    Gf24a4 <= Oc7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Eiwla4 <= 1'b1;
	end
	else
	  begin
	    Eiwla4 <= Eb7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ekwla4 <= 1'b1;
	end
	else
	  begin
	    Ekwla4 <= U97x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Emwla4 <= 1'b1;
	end
	else
	  begin
	    Emwla4 <= Ke7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Dowla4 <= 1'b1;
	end
	else
	  begin
	    Dowla4 <= Ag4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cqwla4 <= 1'b0;
	end
	else
	  begin
	    Cqwla4 <= A74x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Dswla4 <= 1'b1;
	end
	else
	  begin
	    Dswla4 <= Qe7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cuwla4 <= 1'b1;
	end
	else
	  begin
	    Cuwla4 <= Ee7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Bwwla4 <= 1'b1;
	end
	else
	  begin
	    Bwwla4 <= Ou7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Aywla4 <= 1'b1;
	end
	else
	  begin
	    Aywla4 <= Mp6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Zzwla4 <= 1'b1;
	end
	else
	  begin
	    Zzwla4 <= Kn5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Z1xla4 <= 1'b1;
	end
	else
	  begin
	    Z1xla4 <= Qn5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Z3xla4 <= 1'b1;
	end
	else
	  begin
	    Z3xla4 <= Wn5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Z5xla4 <= 1'b1;
	end
	else
	  begin
	    Z5xla4 <= Co5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Z7xla4 <= 1'b1;
	end
	else
	  begin
	    Z7xla4 <= Io5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Z9xla4 <= 1'b1;
	end
	else
	  begin
	    Z9xla4 <= Oo5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Zbxla4 <= 1'b1;
	end
	else
	  begin
	    Zbxla4 <= Ap5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Zdxla4 <= 1'b1;
	end
	else
	  begin
	    Zdxla4 <= Mp5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Zfxla4 <= 1'b1;
	end
	else
	  begin
	    Zfxla4 <= Sp5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Zhxla4 <= 1'b1;
	end
	else
	  begin
	    Zhxla4 <= Yp5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Zjxla4 <= 1'b1;
	end
	else
	  begin
	    Zjxla4 <= Eq5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Zlxla4 <= 1'b1;
	end
	else
	  begin
	    Zlxla4 <= Kq5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Znxla4 <= 1'b1;
	end
	else
	  begin
	    Znxla4 <= Qq5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Zpxla4 <= 1'b1;
	end
	else
	  begin
	    Zpxla4 <= Gp5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Zrxla4 <= 1'b1;
	end
	else
	  begin
	    Zrxla4 <= Uo5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ztxla4 <= 1'b1;
	end
	else
	  begin
	    Ztxla4 <= En5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Zvxla4 <= 1'b1;
	end
	else
	  begin
	    Zvxla4 <= Ms7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Yxxla4 <= 1'b1;
	end
	else
	  begin
	    Yxxla4 <= Q56x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Yzxla4 <= 1'b1;
	end
	else
	  begin
	    Yzxla4 <= W56x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Y1yla4 <= 1'b1;
	end
	else
	  begin
	    Y1yla4 <= C66x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Y3yla4 <= 1'b1;
	end
	else
	  begin
	    Y3yla4 <= I66x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Y5yla4 <= 1'b1;
	end
	else
	  begin
	    Y5yla4 <= O66x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Y7yla4 <= 1'b1;
	end
	else
	  begin
	    Y7yla4 <= U66x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Y9yla4 <= 1'b1;
	end
	else
	  begin
	    Y9yla4 <= A76x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ybyla4 <= 1'b1;
	end
	else
	  begin
	    Ybyla4 <= G76x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ydyla4 <= 1'b1;
	end
	else
	  begin
	    Ydyla4 <= M76x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Yfyla4 <= 1'b1;
	end
	else
	  begin
	    Yfyla4 <= S76x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Yhyla4 <= 1'b1;
	end
	else
	  begin
	    Yhyla4 <= Y76x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Yjyla4 <= 1'b1;
	end
	else
	  begin
	    Yjyla4 <= E86x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ylyla4 <= 1'b1;
	end
	else
	  begin
	    Ylyla4 <= K86x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ynyla4 <= 1'b1;
	end
	else
	  begin
	    Ynyla4 <= Q86x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ypyla4 <= 1'b1;
	end
	else
	  begin
	    Ypyla4 <= W86x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Yryla4 <= 1'b1;
	end
	else
	  begin
	    Yryla4 <= C96x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ytyla4 <= 1'b1;
	end
	else
	  begin
	    Ytyla4 <= Ss7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xvyla4 <= 1'b1;
	end
	else
	  begin
	    Xvyla4 <= O97x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xxyla4 <= 1'b1;
	end
	else
	  begin
	    Xxyla4 <= Ya7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xzyla4 <= 1'b1;
	end
	else
	  begin
	    Xzyla4 <= Ic7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  X1zla4 <= 1'b1;
	end
	else
	  begin
	    X1zla4 <= Sd7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  X3zla4 <= 1'b1;
	end
	else
	  begin
	    X3zla4 <= Cf7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  X5zla4 <= 1'b1;
	end
	else
	  begin
	    X5zla4 <= Mg7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  X7zla4 <= 1'b1;
	end
	else
	  begin
	    X7zla4 <= Sj7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  X9zla4 <= 1'b1;
	end
	else
	  begin
	    X9zla4 <= Mm7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xbzla4 <= 1'b1;
	end
	else
	  begin
	    Xbzla4 <= Gp7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xdzla4 <= 1'b1;
	end
	else
	  begin
	    Xdzla4 <= Qq7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xfzla4 <= 1'b1;
	end
	else
	  begin
	    Xfzla4 <= Am8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xhzla4 <= 1'b1;
	end
	else
	  begin
	    Xhzla4 <= Wn7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xjzla4 <= 1'b1;
	end
	else
	  begin
	    Xjzla4 <= Cl7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xlzla4 <= 1'b1;
	end
	else
	  begin
	    Xlzla4 <= Aj7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xnzla4 <= 1'b1;
	end
	else
	  begin
	    Xnzla4 <= Ci7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xpzla4 <= 1'b1;
	end
	else
	  begin
	    Xpzla4 <= Oo4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xrzla4 <= 1'b1;
	end
	else
	  begin
	    Xrzla4 <= Ys7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Wtzla4 <= 1'b1;
	end
	else
	  begin
	    Wtzla4 <= E58x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Vvzla4 <= 1'b0;
	end
	else
	  begin
	    Vvzla4 <= O98x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Uxzla4 <= 1'b1;
	end
	else
	  begin
	    Uxzla4 <= Ucax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Vzzla4 <= 1'b1;
	end
	else
	  begin
	    Vzzla4 <= Pdax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  W10ma4 <= 1'b1;
	end
	else
	  begin
	    W10ma4 <= A17x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  T30ma4 <= 1'b1;
	end
	else
	  begin
	    T30ma4 <= Dlax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  T50ma4 <= 1'b1;
	end
	else
	  begin
	    T50ma4 <= Sj5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  T70ma4 <= 1'b1;
	end
	else
	  begin
	    T70ma4 <= Yj5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  T90ma4 <= 1'b1;
	end
	else
	  begin
	    T90ma4 <= Ek5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Tb0ma4 <= 1'b1;
	end
	else
	  begin
	    Tb0ma4 <= Kk5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Td0ma4 <= 1'b1;
	end
	else
	  begin
	    Td0ma4 <= Qk5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Tf0ma4 <= 1'b1;
	end
	else
	  begin
	    Tf0ma4 <= Wk5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Th0ma4 <= 1'b1;
	end
	else
	  begin
	    Th0ma4 <= Il5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Tj0ma4 <= 1'b1;
	end
	else
	  begin
	    Tj0ma4 <= Ul5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Tl0ma4 <= 1'b1;
	end
	else
	  begin
	    Tl0ma4 <= Am5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Tn0ma4 <= 1'b1;
	end
	else
	  begin
	    Tn0ma4 <= Gm5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Tp0ma4 <= 1'b1;
	end
	else
	  begin
	    Tp0ma4 <= Mm5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Tr0ma4 <= 1'b1;
	end
	else
	  begin
	    Tr0ma4 <= Sm5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Tt0ma4 <= 1'b1;
	end
	else
	  begin
	    Tt0ma4 <= Ym5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Tv0ma4 <= 1'b1;
	end
	else
	  begin
	    Tv0ma4 <= Ol5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Tx0ma4 <= 1'b1;
	end
	else
	  begin
	    Tx0ma4 <= Cl5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Tz0ma4 <= 1'b1;
	end
	else
	  begin
	    Tz0ma4 <= Mj5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  T11ma4 <= 1'b1;
	end
	else
	  begin
	    T11ma4 <= Kz7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Q31ma4 <= 1'b1;
	end
	else
	  begin
	    Q31ma4 <= Tmax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Q51ma4 <= 1'b1;
	end
	else
	  begin
	    Q51ma4 <= Y16x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Q71ma4 <= 1'b1;
	end
	else
	  begin
	    Q71ma4 <= O36x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Q91ma4 <= 1'b1;
	end
	else
	  begin
	    Q91ma4 <= A46x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Qb1ma4 <= 1'b1;
	end
	else
	  begin
	    Qb1ma4 <= K56x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Qd1ma4 <= 1'b1;
	end
	else
	  begin
	    Qd1ma4 <= E56x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Qf1ma4 <= 1'b1;
	end
	else
	  begin
	    Qf1ma4 <= Y46x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Qh1ma4 <= 1'b1;
	end
	else
	  begin
	    Qh1ma4 <= S46x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Qj1ma4 <= 1'b1;
	end
	else
	  begin
	    Qj1ma4 <= M46x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ql1ma4 <= 1'b1;
	end
	else
	  begin
	    Ql1ma4 <= G46x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Qn1ma4 <= 1'b1;
	end
	else
	  begin
	    Qn1ma4 <= U36x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Qp1ma4 <= 1'b1;
	end
	else
	  begin
	    Qp1ma4 <= I36x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Qr1ma4 <= 1'b1;
	end
	else
	  begin
	    Qr1ma4 <= C36x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Qt1ma4 <= 1'b1;
	end
	else
	  begin
	    Qt1ma4 <= W26x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Qv1ma4 <= 1'b1;
	end
	else
	  begin
	    Qv1ma4 <= Q26x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Qx1ma4 <= 1'b1;
	end
	else
	  begin
	    Qx1ma4 <= K26x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Qz1ma4 <= 1'b1;
	end
	else
	  begin
	    Qz1ma4 <= E26x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Q12ma4 <= 1'b1;
	end
	else
	  begin
	    Q12ma4 <= Io8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  M32ma4 <= 1'b1;
	end
	else
	  begin
	    M32ma4 <= Vnax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  L52ma4 <= 1'b1;
	end
	else
	  begin
	    L52ma4 <= Sg6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  K72ma4 <= 1'b1;
	end
	else
	  begin
	    K72ma4 <= Yg6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  J92ma4 <= 1'b1;
	end
	else
	  begin
	    J92ma4 <= Eh6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ib2ma4 <= 1'b1;
	end
	else
	  begin
	    Ib2ma4 <= Kh6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hd2ma4 <= 1'b1;
	end
	else
	  begin
	    Hd2ma4 <= Qh6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Gf2ma4 <= 1'b1;
	end
	else
	  begin
	    Gf2ma4 <= Wh6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Fh2ma4 <= 1'b1;
	end
	else
	  begin
	    Fh2ma4 <= Ci6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ej2ma4 <= 1'b1;
	end
	else
	  begin
	    Ej2ma4 <= Ii6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Dl2ma4 <= 1'b1;
	end
	else
	  begin
	    Dl2ma4 <= Oi6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cn2ma4 <= 1'b1;
	end
	else
	  begin
	    Cn2ma4 <= Ui6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Bp2ma4 <= 1'b1;
	end
	else
	  begin
	    Bp2ma4 <= Aj6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ar2ma4 <= 1'b1;
	end
	else
	  begin
	    Ar2ma4 <= Gj6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Zs2ma4 <= 1'b1;
	end
	else
	  begin
	    Zs2ma4 <= Mj6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Yu2ma4 <= 1'b1;
	end
	else
	  begin
	    Yu2ma4 <= Sj6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xw2ma4 <= 1'b1;
	end
	else
	  begin
	    Xw2ma4 <= Yj6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Wy2ma4 <= 1'b1;
	end
	else
	  begin
	    Wy2ma4 <= Ek6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  V03ma4 <= 1'b1;
	end
	else
	  begin
	    V03ma4 <= Qk6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  U23ma4 <= 1'b1;
	end
	else
	  begin
	    U23ma4 <= Wk6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  T43ma4 <= 1'b1;
	end
	else
	  begin
	    T43ma4 <= Cl6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  S63ma4 <= 1'b1;
	end
	else
	  begin
	    S63ma4 <= Il6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  R83ma4 <= 1'b1;
	end
	else
	  begin
	    R83ma4 <= Ol6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Qa3ma4 <= 1'b1;
	end
	else
	  begin
	    Qa3ma4 <= Ul6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Pc3ma4 <= 1'b1;
	end
	else
	  begin
	    Pc3ma4 <= Gm6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Oe3ma4 <= 1'b1;
	end
	else
	  begin
	    Oe3ma4 <= Sm6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ng3ma4 <= 1'b1;
	end
	else
	  begin
	    Ng3ma4 <= Ym6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mi3ma4 <= 1'b1;
	end
	else
	  begin
	    Mi3ma4 <= En6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Lk3ma4 <= 1'b1;
	end
	else
	  begin
	    Lk3ma4 <= Kn6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Km3ma4 <= 1'b1;
	end
	else
	  begin
	    Km3ma4 <= Qn6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Jo3ma4 <= 1'b1;
	end
	else
	  begin
	    Jo3ma4 <= Wn6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Iq3ma4 <= 1'b1;
	end
	else
	  begin
	    Iq3ma4 <= Mm6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hs3ma4 <= 1'b1;
	end
	else
	  begin
	    Hs3ma4 <= Am6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Gu3ma4 <= 1'b1;
	end
	else
	  begin
	    Gu3ma4 <= Kk6x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Fw3ma4 <= 1'b1;
	end
	else
	  begin
	    Fw3ma4 <= Ez7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cy3ma4 <= 1'b0;
	end
	else
	  begin
	    Cy3ma4 <= Yj8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  D04ma4 <= 1'b0;
	end
	else
	  begin
	    D04ma4 <= Sj8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  E24ma4 <= 1'b0;
	end
	else
	  begin
	    E24ma4 <= Ek8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  F44ma4 <= 1'b0;
	end
	else
	  begin
	    F44ma4 <= W88x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  E64ma4 <= 1'b0;
	end
	else
	  begin
	    E64ma4 <= C98x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  D84ma4 <= 1'b0;
	end
	else
	  begin
	    D84ma4 <= U08x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Fa4ma4 <= 1'b0;
	end
	else
	  begin
	    Fa4ma4 <= G18x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hc4ma4 <= 1'b0;
	end
	else
	  begin
	    Hc4ma4 <= Wz7x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Je4ma4 <= 1'b0;
	end
	else
	  begin
	    Je4ma4 <= Qn8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Lg4ma4 <= 1'b0;
	end
	else
	  begin
	    Lg4ma4 <= Kh8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ni4ma4 <= 1'b0;
	end
	else
	  begin
	    Ni4ma4 <= Qh8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Pk4ma4 <= 1'b0;
	end
	else
	  begin
	    Pk4ma4 <= Eh8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Qm4ma4 <= 1'b0;
	end
	else
	  begin
	    Qm4ma4 <= Ga8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ro4ma4 <= 1'b0;
	end
	else
	  begin
	    Ro4ma4 <= Aa8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Sq4ma4 <= 1'b0;
	end
	else
	  begin
	    Sq4ma4 <= I98x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ss4ma4 <= 1'b0;
	end
	else
	  begin
	    Ss4ma4 <= Ye63a4;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Uu4ma4 <= 1'b0;
	end
	else
	  begin
	    Uu4ma4 <= Ff63a4;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ww4ma4 <= 1'b0;
	end
	else
	  begin
	    Ww4ma4 <= Re63a4;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Yy4ma4 <= 1'b0;
	end
	else
	  begin
	    Yy4ma4 <= Mf63a4;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  A15ma4 <= 1'b0;
	end
	else
	  begin
	    A15ma4 <= Wh8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  A35ma4 <= 1'b0;
	end
	else
	  begin
	    A35ma4 <= Ci8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  A55ma4 <= 1'b0;
	end
	else
	  begin
	    A55ma4 <= Ii8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  A75ma4 <= 1'b0;
	end
	else
	  begin
	    A75ma4 <= Mj8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  A95ma4 <= 1'b1;
	end
	else
	  begin
	    A95ma4 <= If8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Cb5ma4 <= 1'b1;
	end
	else
	  begin
	    Cb5ma4 <= Vgax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ed5ma4 <= 1'b1;
	end
	else
	  begin
	    Ed5ma4 <= Yd8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ff5ma4 <= 1'b1;
	end
	else
	  begin
	    Ff5ma4 <= Ffax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Gh5ma4 <= 1'b1;
	end
	else
	  begin
	    Gh5ma4 <= Md8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hj5ma4 <= 1'b1;
	end
	else
	  begin
	    Hj5ma4 <= Reax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Il5ma4 <= 1'b1;
	end
	else
	  begin
	    Il5ma4 <= Gd8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Jn5ma4 <= 1'b1;
	end
	else
	  begin
	    Jn5ma4 <= Keax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Kp5ma4 <= 1'b1;
	end
	else
	  begin
	    Kp5ma4 <= Ad8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Lr5ma4 <= 1'b1;
	end
	else
	  begin
	    Lr5ma4 <= Deax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Mt5ma4 <= 1'b1;
	end
	else
	  begin
	    Mt5ma4 <= Uc8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Nv5ma4 <= 1'b1;
	end
	else
	  begin
	    Nv5ma4 <= Wdax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ox5ma4 <= 1'b1;
	end
	else
	  begin
	    Ox5ma4 <= Oc8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Pz5ma4 <= 1'b1;
	end
	else
	  begin
	    Pz5ma4 <= Ic8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Q16ma4 <= 1'b1;
	end
	else
	  begin
	    Q16ma4 <= Cc8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  R36ma4 <= 1'b1;
	end
	else
	  begin
	    R36ma4 <= Wb8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  S56ma4 <= 1'b1;
	end
	else
	  begin
	    S56ma4 <= Coax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  R76ma4 <= 1'b1;
	end
	else
	  begin
	    R76ma4 <= Yj4x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  R96ma4 <= 1'b1;
	end
	else
	  begin
	    R96ma4 <= Pkax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rb6ma4 <= 1'b1;
	end
	else
	  begin
	    Rb6ma4 <= Cc5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rd6ma4 <= 1'b1;
	end
	else
	  begin
	    Rd6ma4 <= Sd5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rf6ma4 <= 1'b1;
	end
	else
	  begin
	    Rf6ma4 <= Ee5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rh6ma4 <= 1'b1;
	end
	else
	  begin
	    Rh6ma4 <= Of5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rj6ma4 <= 1'b1;
	end
	else
	  begin
	    Rj6ma4 <= If5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rl6ma4 <= 1'b1;
	end
	else
	  begin
	    Rl6ma4 <= Cf5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rn6ma4 <= 1'b1;
	end
	else
	  begin
	    Rn6ma4 <= We5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rp6ma4 <= 1'b1;
	end
	else
	  begin
	    Rp6ma4 <= Qe5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rr6ma4 <= 1'b1;
	end
	else
	  begin
	    Rr6ma4 <= Ke5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rt6ma4 <= 1'b1;
	end
	else
	  begin
	    Rt6ma4 <= Yd5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rv6ma4 <= 1'b1;
	end
	else
	  begin
	    Rv6ma4 <= Md5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rx6ma4 <= 1'b1;
	end
	else
	  begin
	    Rx6ma4 <= Gd5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Rz6ma4 <= 1'b1;
	end
	else
	  begin
	    Rz6ma4 <= Ad5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  R17ma4 <= 1'b1;
	end
	else
	  begin
	    R17ma4 <= Uc5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  R37ma4 <= 1'b1;
	end
	else
	  begin
	    R37ma4 <= Oc5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  R57ma4 <= 1'b1;
	end
	else
	  begin
	    R57ma4 <= Ic5x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  R77ma4 <= 1'b1;
	end
	else
	  begin
	    R77ma4 <= Sg8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  T97ma4 <= 1'b1;
	end
	else
	  begin
	    T97ma4 <= Liax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Vb7ma4 <= 1'b1;
	end
	else
	  begin
	    Vb7ma4 <= Sd8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Wd7ma4 <= 1'b1;
	end
	else
	  begin
	    Wd7ma4 <= Yeax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Xf7ma4 <= 1'b1;
	end
	else
	  begin
	    Xf7ma4 <= We8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Zh7ma4 <= 1'b1;
	end
	else
	  begin
	    Zh7ma4 <= Hgax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Bk7ma4 <= 1'b1;
	end
	else
	  begin
	    Bk7ma4 <= Gg8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Dm7ma4 <= 1'b1;
	end
	else
	  begin
	    Dm7ma4 <= Xhax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Fo7ma4 <= 1'b1;
	end
	else
	  begin
	    Fo7ma4 <= Idax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Gq7ma4 <= 1'b1;
	end
	else
	  begin
	    Gq7ma4 <= Bdax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hs7ma4 <= 1'b0;
	end
	else
	  begin
	    Hs7ma4 <= U64x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Iu7ma4 <= 1'b0;
	end
	else
	  begin
	    Iu7ma4 <= K88x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Hw7ma4 <= 1'b1;
	end
	else
	  begin
	    Hw7ma4 <= Yg8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Jy7ma4 <= 1'b1;
	end
	else
	  begin
	    Jy7ma4 <= Siax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  L08ma4 <= 1'b0;
	end
	else
	  begin
	    L08ma4 <= Sa8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  M28ma4 <= 1'b1;
	end
	else
	  begin
	    M28ma4 <= Kq8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  O48ma4 <= 1'b0;
	end
	else
	  begin
	    O48ma4 <= Ma8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  P68ma4 <= 1'b1;
	end
	else
	  begin
	    P68ma4 <= Cf8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  R88ma4 <= 1'b1;
	end
	else
	  begin
	    R88ma4 <= Ogax84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ta8ma4 <= 1'b0;
	end
	else
	  begin
	    Ta8ma4 <= Eb8x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Uc8ma4 <= 1'b0;
	end
	else
	  begin
	    Uc8ma4 <= O64x84;
	  end
	always @(posedge HCLK or negedge HRESETn) if (~HRESETn) begin
	  Ve8ma4 <= 1'b0;
	end
	else
	  begin
	    Ve8ma4 <= I64x84;
	  end
endmodule

// ===================
//  DESIGN STATISTICS 
// ===================
//                                        Static<!>  Elaborated<@>
//                                        ------     ----------
// No. of module instances:                    1              1
// No. of comb. udp instances:                 0              0
// No. of seq. udp instances:                  0              0
// No. of gates:                               0              0
// No. of (r)tran(if[01])s:                    0              0
// No. of continuous assignments:          10487          10487
// No. of module+udp port connects:            0              0
// No. of registers (vector+scalar):         783            783
// No. of memories:                            0              0
// No. of scalar nets:                     10335          10335
// No. of vector nets:                        27             27
// No. of named events:                        0              0
// No. of always blocks:                     783            783
// No. of initial blocks:                      0              0
// No. of fork/join blocks:                    0              0
// No. of verilog tasks:                       0              0
// No. of verilog functions:                   0              0
// No. of verilog task calls:                  0              0
// No. of verilog function calls:              0              0
// No. of system task calls:                   0              0
// No. of user task calls:                     0              0
// No. of system function calls:               0              0
// No. of user function calls:                 0              0
// No. of hierarchical references:             0              0
// No. of concatenations:                     13             13
// No. of force/release statements:            0              0
// No. of bit selects:                      1094           1094
// No. of part selects:                        4              4
// No. of non-blocking assignments:         1566           1566
// No. of specify blocks<#>:                   0              0
// No. of timing checks:                       0              0
//
// No. of top level modules:                   1
//        modules:                             1
// No. of udps:                                0
//        seq. udps:                           0
//        comb. udps:                          0
// No. of module+udp ports:                   25
// No. of system tasks:                        0
// No. of user tasks:                          0
// No. of system functions:                    0
// No. of user functions:                      0
//
// Footnotes:
// ---------
// <!> No. of unique instances of a construct as it appears in the source.
// <@> No. of instances of a construct when the design is elaborated.
// <#> Multiple specify blocks in the SAME module are combined and counted
//     as ONE block.
